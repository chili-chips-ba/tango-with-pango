//
// Generated (version 2022.2-SP4.2<build 132111>) at Mon Oct 23 14:00:24 2023
//

module top_lcd_touch
(
    input sys_clk,
    input sys_rst_n,
    output lcd_bl,
    output lcd_clk,
    output lcd_de,
    output lcd_hs,
    output lcd_rst_n,
    output lcd_vs,
    output touch_rst_n,
    output touch_scl,
    inout [23:0] lcd_rgb,
    inout touch_int,
    inout touch_sda
);
	// SDC constraint : (object sys_clk) (id 1000) (clock sys_clk) (249 : D:/Desktop/50G/29_top_lcd_touch/prj/top_lcd_touch.fdc)
    wire _N0;
    wire _N1;
    wire _N2;
    wire _N3;
    wire _N48;
    wire _N68;
    wire _N88;
    wire _N108;
    wire _N154;
    wire _N174;
    wire _N194;
    wire _N574;
    wire _N619;
    wire _N620;
    wire _N621;
    wire _N622;
    wire _N623;
    wire _N624;
    wire _N625;
    wire _N627;
    wire _N628;
    wire _N629;
    wire _N630;
    wire _N631;
    wire _N632;
    wire _N633;
    wire _N634;
    wire _N636;
    wire _N637;
    wire _N638;
    wire _N639;
    wire _N640;
    wire _N641;
    wire _N642;
    wire _N643;
    wire _N645;
    wire _N646;
    wire _N647;
    wire _N648;
    wire _N649;
    wire _N650;
    wire _N651;
    wire _N652;
    wire _N653;
    wire _N655;
    wire _N656;
    wire _N657;
    wire _N658;
    wire _N659;
    wire _N660;
    wire _N661;
    wire _N662;
    wire _N663;
    wire _N664;
    wire _N665;
    wire _N666;
    wire _N667;
    wire _N668;
    wire _N669;
    wire _N670;
    wire _N671;
    wire _N672;
    wire _N673;
    wire _N675;
    wire _N676;
    wire _N677;
    wire _N678;
    wire _N679;
    wire _N680;
    wire _N682;
    wire _N683;
    wire _N684;
    wire _N685;
    wire _N686;
    wire _N687;
    wire _N688;
    wire _N690;
    wire _N691;
    wire _N692;
    wire _N693;
    wire _N694;
    wire _N695;
    wire _N696;
    wire _N697;
    wire _N698;
    wire _N700;
    wire _N701;
    wire _N702;
    wire _N703;
    wire _N704;
    wire _N705;
    wire _N706;
    wire _N707;
    wire _N708;
    wire _N709;
    wire _N711;
    wire _N712;
    wire _N713;
    wire _N714;
    wire _N715;
    wire _N716;
    wire _N717;
    wire _N718;
    wire _N719;
    wire _N720;
    wire _N722;
    wire _N723;
    wire _N724;
    wire _N725;
    wire _N726;
    wire _N728;
    wire _N729;
    wire _N730;
    wire _N731;
    wire _N784;
    wire _N785;
    wire _N791;
    wire _N2517;
    wire _N2521;
    wire _N2528;
    wire _N2543;
    wire _N2552;
    wire _N2555;
    wire _N2558;
    wire _N2560;
    wire _N2571;
    wire _N2574;
    wire _N2576;
    wire _N2577;
    wire _N2578;
    wire _N4964;
    wire _N5000;
    wire _N5003;
    wire _N5005;
    wire _N5007;
    wire _N9388;
    wire _N9402;
    wire _N9403;
    wire _N9426;
    wire _N9468;
    wire _N9512;
    wire _N9551;
    wire _N9596;
    wire _N9641;
    wire _N9679;
    wire _N9724;
    wire _N9759;
    wire _N9791;
    wire _N9827;
    wire _N9859;
    wire _N9907;
    wire _N9955;
    wire _N10009;
    wire _N10046;
    wire _N10093;
    wire _N10183_5;
    wire _N10183_6;
    wire _N10183_7;
    wire _N10183_9;
    wire _N10183_11;
    wire _N10183_12;
    wire _N10183_17;
    wire _N10183_18;
    wire _N10183_20;
    wire _N10183_21;
    wire _N10183_22;
    wire _N10183_23;
    wire _N10183_24;
    wire _N10183_25;
    wire _N10183_26;
    wire _N10183_28;
    wire _N10183_31;
    wire _N10183_36;
    wire _N10183_40;
    wire _N10183_41;
    wire _N10183_42;
    wire _N10183_43;
    wire _N10183_44;
    wire _N10183_45;
    wire _N10183_46;
    wire _N10183_47;
    wire _N10183_48;
    wire _N10183_49;
    wire _N10183_50;
    wire _N10183_51;
    wire _N10183_52;
    wire _N10183_53;
    wire _N10183_58;
    wire _N10183_59;
    wire _N10183_62;
    wire _N10183_69;
    wire _N10183_71;
    wire _N10183_73;
    wire _N10183_75;
    wire _N10183_77;
    wire _N10183_79;
    wire _N10183_81;
    wire _N10183_83;
    wire _N10183_84;
    wire _N10183_85;
    wire _N10183_86;
    wire _N10183_87_inv;
    wire _N10183_88;
    wire _N10183_89;
    wire _N10183_90;
    wire _N10183_91_inv;
    wire _N10183_92;
    wire _N10183_93;
    wire _N10183_94;
    wire _N10183_95_inv;
    wire _N10183_97;
    wire _N10183_98;
    wire _N10183_101;
    wire _N10183_102;
    wire _N10183_104;
    wire _N10183_105;
    wire _N10183_106;
    wire _N10183_108;
    wire _N10183_109;
    wire _N10183_112;
    wire _N10183_113;
    wire _N10183_114;
    wire _N10183_116;
    wire _N10183_117;
    wire _N10183_120;
    wire _N10183_121;
    wire _N10183_122;
    wire _N10183_124;
    wire _N10183_125;
    wire _N10183_128;
    wire _N10183_129;
    wire _N10183_130;
    wire _N10183_132;
    wire _N10183_133;
    wire _N10183_137;
    wire _N10183_138;
    wire _N10183_140;
    wire _N10183_145;
    wire _N10183_146;
    wire _N10183_148;
    wire _N10183_153;
    wire _N10183_154;
    wire _N10183_156;
    wire _N10183_160;
    wire _N10183_162;
    wire _N10183_163;
    wire _N10183_166;
    wire _N10183_167;
    wire _N10183_168;
    wire _N10183_171;
    wire _N10183_172;
    wire _N10183_174;
    wire _N10183_175;
    wire _N10183_176;
    wire _N10183_177;
    wire _N10183_178;
    wire _N10183_180;
    wire _N10183_181;
    wire _N10183_182;
    wire _N10183_184;
    wire _N10183_185;
    wire _N10183_186;
    wire _N10183_187;
    wire _N10183_188;
    wire _N10183_189;
    wire _N10183_190;
    wire _N10183_191;
    wire _N10183_192;
    wire _N10183_193;
    wire _N10183_194;
    wire _N10183_196;
    wire _N10183_197;
    wire _N10183_198;
    wire _N10183_200;
    wire _N10183_201;
    wire _N10183_202;
    wire _N10183_203;
    wire _N10183_204;
    wire _N10183_205;
    wire _N10183_206;
    wire _N10183_207;
    wire _N10183_208;
    wire _N10183_209;
    wire _N10183_210;
    wire _N10183_212;
    wire _N10183_213;
    wire _N10183_214;
    wire _N10183_216;
    wire _N10183_217;
    wire _N10183_218;
    wire _N10183_219;
    wire _N10183_220;
    wire _N10183_221;
    wire _N10183_222;
    wire _N10183_223;
    wire _N10183_224;
    wire _N10183_225;
    wire _N10183_226;
    wire _N10183_228;
    wire _N10183_229;
    wire _N10183_230;
    wire _N10183_232;
    wire _N10183_233;
    wire _N10183_234;
    wire _N10183_235;
    wire _N10183_236;
    wire _N10183_237;
    wire _N10183_238;
    wire _N10183_239;
    wire _N10183_240;
    wire _N10183_241;
    wire _N10183_242;
    wire _N10183_244;
    wire _N10183_245;
    wire _N10183_246;
    wire _N10183_248;
    wire _N10183_249;
    wire _N10183_250;
    wire _N10183_251;
    wire _N10183_252;
    wire _N10183_253;
    wire _N10183_254;
    wire _N10183_255;
    wire _N10183_256;
    wire _N10183_257;
    wire _N10183_258;
    wire _N10183_260;
    wire _N10183_261;
    wire _N10183_262;
    wire _N10183_264;
    wire _N10183_265;
    wire _N10183_266;
    wire _N10183_267;
    wire _N10183_268;
    wire _N10183_269;
    wire _N10183_270;
    wire _N10183_271;
    wire _N10183_272;
    wire _N10183_273;
    wire _N10183_274;
    wire _N10183_276;
    wire _N10183_277;
    wire _N10183_278;
    wire _N10183_280;
    wire _N10183_281;
    wire _N10183_282;
    wire _N10183_283;
    wire _N10183_284;
    wire _N10183_286;
    wire _N10183_288;
    wire _N10183_290;
    wire _N10183_292;
    wire _N10183_295;
    wire _N10183_296;
    wire _N10183_300;
    wire _N10183_301;
    wire _N10183_302;
    wire _N10183_306;
    wire _N10183_307;
    wire _N10183_309;
    wire _N10183_310;
    wire _N10183_311;
    wire _N10183_312;
    wire _N10183_315;
    wire _N10183_317;
    wire _N10183_318;
    wire _N10183_319_inv;
    wire _N10183_320;
    wire _N10183_321;
    wire _N10183_322;
    wire _N10183_323_inv;
    wire _N10183_324;
    wire _N10183_325;
    wire _N10183_328;
    wire _N10183_330;
    wire _N10183_331_inv;
    wire _N10183_332;
    wire _N10183_333;
    wire _N10183_334;
    wire _N10183_335;
    wire _N10183_336;
    wire _N10183_338;
    wire _N10183_339;
    wire _N10183_341;
    wire _N10183_342;
    wire _N10183_343;
    wire _N10183_344;
    wire _N10183_347;
    wire _N10183_349;
    wire _N10183_350_inv;
    wire _N10183_351;
    wire _N10183_352;
    wire _N10183_353;
    wire _N10183_354_inv;
    wire _N10183_355;
    wire _N10183_356;
    wire _N10183_359;
    wire _N10183_361;
    wire _N10183_362_inv;
    wire _N10183_363;
    wire _N10183_364;
    wire _N10183_365;
    wire _N10183_366;
    wire _N10183_367;
    wire _N10183_369;
    wire _N10183_370;
    wire _N10183_372;
    wire _N10183_373;
    wire _N10183_374;
    wire _N10183_375;
    wire _N10183_378;
    wire _N10183_380;
    wire _N10183_381_inv;
    wire _N10183_382;
    wire _N10183_383;
    wire _N10183_384;
    wire _N10183_385_inv;
    wire _N10183_386;
    wire _N10183_387;
    wire _N10183_390;
    wire _N10183_392;
    wire _N10183_393_inv;
    wire _N10183_394;
    wire _N10183_395;
    wire _N10183_396;
    wire _N10183_397;
    wire _N10183_398;
    wire _N10183_400;
    wire _N10183_401;
    wire _N10183_403;
    wire _N10183_404;
    wire _N10183_405;
    wire _N10183_406;
    wire _N10183_409;
    wire _N10183_411;
    wire _N10183_412_inv;
    wire _N10183_413;
    wire _N10183_414;
    wire _N10183_415;
    wire _N10183_416_inv;
    wire _N10183_417;
    wire _N10183_418;
    wire _N10183_421;
    wire _N10183_423;
    wire _N10183_424_inv;
    wire _N10183_425;
    wire _N10183_426;
    wire _N10183_427;
    wire _N10183_428;
    wire _N10183_429;
    wire _N10183_431;
    wire _N10183_432;
    wire _N10183_434;
    wire _N10183_435;
    wire _N10183_436;
    wire _N10183_437;
    wire _N10183_440;
    wire _N10183_442;
    wire _N10183_443_inv;
    wire _N10183_444;
    wire _N10183_445;
    wire _N10183_446;
    wire _N10183_447_inv;
    wire _N10183_448;
    wire _N10183_449;
    wire _N10183_450;
    wire _N10183_452;
    wire _N10183_454;
    wire _N10183_455_inv;
    wire _N10183_456;
    wire _N10183_457;
    wire _N10183_458;
    wire _N10183_459;
    wire _N10183_460;
    wire _N10183_462;
    wire _N10183_463;
    wire _N10183_465;
    wire _N10183_466;
    wire _N10183_467;
    wire _N10183_468;
    wire _N10183_471;
    wire _N10183_473;
    wire _N10183_474_inv;
    wire _N10183_475;
    wire _N10183_476;
    wire _N10183_477;
    wire _N10183_478_inv;
    wire _N10183_479;
    wire _N10183_480;
    wire _N10183_481;
    wire _N10183_483;
    wire _N10183_485;
    wire _N10183_486_inv;
    wire _N10183_487;
    wire _N10183_488;
    wire _N10183_489;
    wire _N10183_490;
    wire _N10183_491;
    wire _N10183_493;
    wire _N10183_494;
    wire _N10183_496;
    wire _N10183_497;
    wire _N10183_498;
    wire _N10183_499;
    wire _N10183_502;
    wire _N10183_504;
    wire _N10183_505_inv;
    wire _N10183_506;
    wire _N10183_507;
    wire _N10183_508;
    wire _N10183_509_inv;
    wire _N10183_510;
    wire _N10183_511;
    wire _N10183_512;
    wire _N10183_514;
    wire _N10183_516;
    wire _N10183_517_inv;
    wire _N10183_518;
    wire _N10183_519;
    wire _N10183_520;
    wire _N10183_521;
    wire _N10183_522;
    wire _N10183_527;
    wire _N10183_534;
    wire _N10183_535;
    wire _N10183_542;
    wire _N10183_543;
    wire _N10183_544;
    wire _N10183_545;
    wire _N10183_546;
    wire _N10183_547;
    wire _N10183_551;
    wire _N10183_554;
    wire _N10183_555;
    wire _N10183_556;
    wire _N10183_558;
    wire _N10183_559;
    wire _N10183_560;
    wire _N10183_561;
    wire _N10183_562;
    wire _N10183_564;
    wire _N10183_571;
    wire _N10183_572;
    wire _N10183_573;
    wire _N10183_574_inv;
    wire _N10183_575;
    wire _N10183_576;
    wire _N10183_577;
    wire _N10183_578;
    wire _N10183_579;
    wire _N10183_580;
    wire _N10183_586;
    wire _N10183_588;
    wire _N10183_589;
    wire _N10183_595;
    wire _N10183_596;
    wire _N10183_597;
    wire _N10183_598;
    wire _N10183_600;
    wire _N10183_601;
    wire _N10183_602;
    wire _N10183_605;
    wire _N10183_611;
    wire _N10183_613;
    wire _N10183_614;
    wire _N10183_616;
    wire _N10183_617;
    wire _N10183_618;
    wire _N10183_619;
    wire _N10183_620;
    wire _N10183_622;
    wire _N10183_628;
    wire _N10183_629;
    wire _N10183_630;
    wire _N10183_631_inv;
    wire _N10183_632;
    wire _N10183_633;
    wire _N10183_634;
    wire _N10183_635;
    wire _N10183_636;
    wire _N10183_642;
    wire _N10183_644;
    wire _N10183_645;
    wire _N10183_651;
    wire _N10183_652;
    wire _N10183_653;
    wire _N10183_654;
    wire _N10183_656;
    wire _N10183_657;
    wire _N10183_658;
    wire _N10183_661;
    wire _N10183_667;
    wire _N10183_669;
    wire _N10183_670;
    wire _N10183_672;
    wire _N10183_673;
    wire _N10183_674;
    wire _N10183_675;
    wire _N10183_676;
    wire _N10183_678;
    wire _N10183_684;
    wire _N10183_685;
    wire _N10183_686;
    wire _N10183_687_inv;
    wire _N10183_688;
    wire _N10183_689;
    wire _N10183_690;
    wire _N10183_691;
    wire _N10183_692;
    wire _N10183_698;
    wire _N10183_700;
    wire _N10183_701;
    wire _N10183_707;
    wire _N10183_708;
    wire _N10183_709;
    wire _N10183_710;
    wire _N10183_712;
    wire _N10183_713;
    wire _N10183_714;
    wire _N10183_717;
    wire _N10183_723;
    wire _N10183_725;
    wire _N10183_726;
    wire _N10183_728;
    wire _N10183_729;
    wire _N10183_730;
    wire _N10183_731;
    wire _N10183_732;
    wire _N10183_734;
    wire _N10183_740;
    wire _N10183_741;
    wire _N10183_742;
    wire _N10183_743_inv;
    wire _N10183_744;
    wire _N10183_745;
    wire _N10183_746;
    wire _N10183_747;
    wire _N10183_748;
    wire _N10183_754;
    wire _N10183_756;
    wire _N10183_757;
    wire _N10183_763;
    wire _N10183_764;
    wire _N10183_765;
    wire _N10183_766;
    wire _N10183_768;
    wire _N10183_769;
    wire _N10183_770;
    wire _N10183_773;
    wire _N10183_779;
    wire _N10183_781;
    wire _N10183_782;
    wire _N10183_784;
    wire _N10183_785;
    wire _N10183_786;
    wire _N10183_787;
    wire _N10183_788;
    wire _N10183_790;
    wire _N10183_796;
    wire _N10183_797;
    wire _N10183_798;
    wire _N10183_799_inv;
    wire _N10183_800;
    wire _N10183_801;
    wire _N10183_802;
    wire _N10183_803;
    wire _N10183_804;
    wire _N10183_810;
    wire _N10183_812;
    wire _N10183_813;
    wire _N10183_819;
    wire _N10183_820;
    wire _N10183_821;
    wire _N10183_822;
    wire _N10183_824;
    wire _N10183_825;
    wire _N10183_826;
    wire _N10183_829;
    wire _N10183_835;
    wire _N10183_837;
    wire _N10183_838;
    wire _N10183_840;
    wire _N10183_841;
    wire _N10183_842;
    wire _N10183_843;
    wire _N10183_844;
    wire _N10183_846;
    wire _N10183_852;
    wire _N10183_853;
    wire _N10183_854;
    wire _N10183_855_inv;
    wire _N10183_856;
    wire _N10183_857;
    wire _N10183_858;
    wire _N10183_859;
    wire _N10183_860;
    wire _N10183_866;
    wire _N10183_868;
    wire _N10183_869;
    wire _N10183_875;
    wire _N10183_876;
    wire _N10183_877;
    wire _N10183_878;
    wire _N10183_880;
    wire _N10183_881;
    wire _N10183_882;
    wire _N10183_885;
    wire _N10183_891;
    wire _N10183_893;
    wire _N10183_894;
    wire _N10183_896;
    wire _N10183_897;
    wire _N10183_898;
    wire _N10183_899;
    wire _N10183_900;
    wire _N10183_902;
    wire _N10183_908;
    wire _N10183_909;
    wire _N10183_910;
    wire _N10183_911_inv;
    wire _N10183_912;
    wire _N10183_913;
    wire _N10183_914;
    wire _N10183_915;
    wire _N10183_916;
    wire _N10183_922;
    wire _N10183_924;
    wire _N10183_925;
    wire _N10183_931;
    wire _N10183_932;
    wire _N10183_933;
    wire _N10183_934;
    wire _N10183_936;
    wire _N10183_937;
    wire _N10183_938;
    wire _N10183_941;
    wire _N10183_947;
    wire _N10183_953;
    wire _N10183_956;
    wire _N10183_957;
    wire _N10183_962;
    wire _N10183_964;
    wire _N10183_966;
    wire _N10183_969;
    wire _N10183_970;
    wire _N10183_974;
    wire _N10183_975;
    wire _N10183_978;
    wire _N10183_983;
    wire _N10183_984;
    wire _N10183_985_inv;
    wire _N10183_988;
    wire _N10183_990;
    wire _N10183_991;
    wire _N10183_992;
    wire _N10183_993;
    wire _N10183_995;
    wire _N10183_996;
    wire _N10183_999;
    wire _N10183_1000;
    wire _N10183_1001_inv;
    wire _N10183_1004;
    wire _N10183_1005;
    wire _N10183_1008;
    wire _N10183_1011_inv;
    wire _N10183_1012;
    wire _N10183_1015;
    wire _N10183_1020_inv;
    wire _N10183_1021;
    wire _N10183_1022_inv;
    wire _N10183_1023;
    wire _N10183_1024;
    wire _N10183_1026;
    wire _N10183_1028;
    wire _N10183_1029;
    wire _N10183_1030;
    wire _N10183_1031;
    wire _N10183_1033;
    wire _N10183_1036;
    wire _N10183_1037;
    wire _N10183_1039;
    wire _N10183_1040;
    wire _N10183_1042;
    wire _N10183_1043;
    wire _N10183_1044;
    wire _N10183_1048;
    wire _N10183_1049;
    wire _N10183_1050;
    wire _N10183_1051;
    wire _N10183_1052;
    wire _N10183_1056;
    wire _N10183_1057;
    wire _N10183_1058_inv;
    wire _N10183_1059;
    wire _N10183_1060;
    wire _N10183_1061;
    wire _N10183_1062_inv;
    wire _N10183_1063;
    wire _N10183_1064;
    wire _N10183_1066;
    wire _N10183_1067;
    wire _N10183_1069;
    wire _N10183_1076;
    wire _N10183_1077;
    wire _N10183_1078_inv;
    wire _N10183_1079;
    wire _N10183_1080;
    wire _N10183_1081_inv;
    wire _N10183_1084;
    wire _N10183_1086;
    wire _N10183_1087;
    wire _N10183_1088;
    wire _N10183_1089;
    wire _N10183_1091;
    wire _N10183_1092;
    wire _N10183_1095;
    wire _N10183_1096;
    wire _N10183_1097_inv;
    wire _N10183_1100;
    wire _N10183_1102;
    wire _N10183_1104_inv;
    wire _N10183_1105;
    wire _N10183_1108;
    wire _N10183_1113_inv;
    wire _N10183_1114;
    wire _N10183_1115_inv;
    wire _N10183_1116;
    wire _N10183_1117;
    wire _N10183_1119;
    wire _N10183_1121;
    wire _N10183_1122;
    wire _N10183_1123;
    wire _N10183_1126;
    wire _N10183_1129;
    wire _N10183_1130;
    wire _N10183_1132;
    wire _N10183_1133;
    wire _N10183_1135;
    wire _N10183_1136;
    wire _N10183_1137;
    wire _N10183_1141;
    wire _N10183_1142;
    wire _N10183_1143;
    wire _N10183_1144;
    wire _N10183_1145;
    wire _N10183_1148;
    wire _N10183_1149;
    wire _N10183_1150_inv;
    wire _N10183_1151;
    wire _N10183_1152;
    wire _N10183_1153;
    wire _N10183_1154_inv;
    wire _N10183_1155;
    wire _N10183_1157;
    wire _N10183_1158;
    wire _N10183_1160;
    wire _N10183_1167;
    wire _N10183_1168;
    wire _N10183_1169_inv;
    wire _N10183_1170;
    wire _N10183_1171;
    wire _N10183_1172_inv;
    wire _N10183_1175;
    wire _N10183_1177;
    wire _N10183_1178;
    wire _N10183_1179;
    wire _N10183_1180;
    wire _N10183_1182;
    wire _N10183_1183;
    wire _N10183_1186;
    wire _N10183_1187;
    wire _N10183_1188_inv;
    wire _N10183_1191;
    wire _N10183_1193;
    wire _N10183_1195_inv;
    wire _N10183_1196;
    wire _N10183_1199;
    wire _N10183_1204_inv;
    wire _N10183_1205;
    wire _N10183_1206_inv;
    wire _N10183_1207;
    wire _N10183_1208;
    wire _N10183_1210;
    wire _N10183_1212;
    wire _N10183_1213;
    wire _N10183_1214;
    wire _N10183_1215;
    wire _N10183_1217;
    wire _N10183_1220;
    wire _N10183_1221;
    wire _N10183_1223;
    wire _N10183_1224;
    wire _N10183_1226;
    wire _N10183_1227;
    wire _N10183_1228;
    wire _N10183_1232;
    wire _N10183_1233;
    wire _N10183_1234;
    wire _N10183_1235;
    wire _N10183_1236;
    wire _N10183_1239;
    wire _N10183_1240;
    wire _N10183_1241_inv;
    wire _N10183_1242;
    wire _N10183_1243;
    wire _N10183_1244;
    wire _N10183_1245_inv;
    wire _N10183_1246;
    wire _N10183_1248;
    wire _N10183_1249;
    wire _N10183_1251;
    wire _N10183_1258;
    wire _N10183_1259;
    wire _N10183_1260_inv;
    wire _N10183_1261;
    wire _N10183_1262;
    wire _N10183_1263_inv;
    wire _N10183_1266;
    wire _N10183_1268;
    wire _N10183_1269;
    wire _N10183_1270;
    wire _N10183_1271;
    wire _N10183_1273;
    wire _N10183_1274;
    wire _N10183_1277;
    wire _N10183_1278;
    wire _N10183_1279_inv;
    wire _N10183_1282;
    wire _N10183_1284;
    wire _N10183_1286_inv;
    wire _N10183_1287;
    wire _N10183_1290;
    wire _N10183_1295_inv;
    wire _N10183_1296;
    wire _N10183_1297_inv;
    wire _N10183_1298;
    wire _N10183_1299;
    wire _N10183_1301;
    wire _N10183_1303;
    wire _N10183_1304;
    wire _N10183_1305;
    wire _N10183_1308;
    wire _N10183_1311;
    wire _N10183_1312;
    wire _N10183_1314;
    wire _N10183_1315;
    wire _N10183_1317;
    wire _N10183_1318;
    wire _N10183_1319;
    wire _N10183_1323;
    wire _N10183_1324;
    wire _N10183_1325;
    wire _N10183_1326;
    wire _N10183_1327;
    wire _N10183_1330;
    wire _N10183_1331;
    wire _N10183_1332_inv;
    wire _N10183_1333;
    wire _N10183_1334;
    wire _N10183_1335;
    wire _N10183_1336_inv;
    wire _N10183_1337;
    wire _N10183_1339;
    wire _N10183_1340;
    wire _N10183_1342;
    wire _N10183_1349;
    wire _N10183_1350;
    wire _N10183_1351_inv;
    wire _N10183_1352;
    wire _N10183_1353;
    wire _N10183_1354_inv;
    wire _N10183_1357;
    wire _N10183_1359;
    wire _N10183_1360;
    wire _N10183_1361;
    wire _N10183_1362;
    wire _N10183_1364;
    wire _N10183_1365;
    wire _N10183_1368;
    wire _N10183_1369;
    wire _N10183_1370_inv;
    wire _N10183_1373;
    wire _N10183_1375;
    wire _N10183_1377_inv;
    wire _N10183_1378;
    wire _N10183_1381;
    wire _N10183_1386_inv;
    wire _N10183_1387;
    wire _N10183_1388_inv;
    wire _N10183_1389;
    wire _N10183_1390;
    wire _N10183_1392;
    wire _N10183_1394;
    wire _N10183_1395;
    wire _N10183_1396;
    wire _N10183_1397;
    wire _N10183_1399;
    wire _N10183_1402;
    wire _N10183_1403;
    wire _N10183_1405;
    wire _N10183_1406;
    wire _N10183_1408;
    wire _N10183_1409;
    wire _N10183_1410;
    wire _N10183_1414;
    wire _N10183_1415;
    wire _N10183_1416;
    wire _N10183_1417;
    wire _N10183_1418;
    wire _N10183_1421;
    wire _N10183_1422;
    wire _N10183_1423_inv;
    wire _N10183_1424;
    wire _N10183_1425;
    wire _N10183_1426;
    wire _N10183_1427_inv;
    wire _N10183_1428;
    wire _N10183_1430;
    wire _N10183_1431;
    wire _N10183_1433;
    wire _N10183_1440;
    wire _N10183_1441;
    wire _N10183_1442_inv;
    wire _N10183_1443;
    wire _N10183_1444;
    wire _N10183_1445_inv;
    wire _N10183_1448;
    wire _N10183_1450;
    wire _N10183_1451;
    wire _N10183_1452;
    wire _N10183_1453;
    wire _N10183_1455;
    wire _N10183_1456;
    wire _N10183_1459;
    wire _N10183_1460;
    wire _N10183_1461_inv;
    wire _N10183_1464;
    wire _N10183_1466;
    wire _N10183_1468_inv;
    wire _N10183_1469;
    wire _N10183_1472;
    wire _N10183_1477_inv;
    wire _N10183_1478;
    wire _N10183_1479_inv;
    wire _N10183_1480;
    wire _N10183_1481;
    wire _N10183_1483;
    wire _N10183_1485;
    wire _N10183_1486;
    wire _N10183_1487;
    wire _N10183_1488;
    wire _N10183_1490;
    wire _N10183_1493;
    wire _N10183_1494;
    wire _N10183_1496;
    wire _N10183_1497;
    wire _N10183_1499;
    wire _N10183_1500;
    wire _N10183_1501;
    wire _N10183_1505;
    wire _N10183_1506;
    wire _N10183_1507;
    wire _N10183_1508;
    wire _N10183_1509;
    wire _N10183_1512;
    wire _N10183_1513;
    wire _N10183_1514_inv;
    wire _N10183_1515;
    wire _N10183_1516;
    wire _N10183_1517;
    wire _N10183_1518_inv;
    wire _N10183_1519;
    wire _N10183_1521;
    wire _N10183_1522;
    wire _N10183_1524;
    wire _N10183_1531;
    wire _N10183_1532;
    wire _N10183_1533_inv;
    wire _N10183_1534;
    wire _N10183_1535;
    wire _N10183_1536_inv;
    wire _N10183_1539;
    wire _N10183_1541;
    wire _N10183_1542;
    wire _N10183_1543;
    wire _N10183_1544;
    wire _N10183_1546;
    wire _N10183_1547;
    wire _N10183_1550;
    wire _N10183_1551;
    wire _N10183_1552_inv;
    wire _N10183_1555;
    wire _N10183_1557;
    wire _N10183_1559_inv;
    wire _N10183_1560;
    wire _N10183_1561;
    wire _N10183_1563;
    wire _N10183_1568_inv;
    wire _N10183_1569;
    wire _N10183_1570_inv;
    wire _N10183_1571;
    wire _N10183_1572;
    wire _N10183_1574;
    wire _N10183_1576;
    wire _N10183_1577;
    wire _N10183_1578;
    wire _N10183_1579;
    wire _N10183_1581;
    wire _N10183_1584;
    wire _N10183_1585;
    wire _N10183_1587;
    wire _N10183_1588;
    wire _N10183_1590;
    wire _N10183_1591;
    wire _N10183_1592;
    wire _N10183_1596;
    wire _N10183_1597;
    wire _N10183_1598;
    wire _N10183_1599;
    wire _N10183_1600;
    wire _N10183_1603;
    wire _N10183_1604;
    wire _N10183_1605_inv;
    wire _N10183_1606;
    wire _N10183_1607;
    wire _N10183_1608;
    wire _N10183_1609_inv;
    wire _N10183_1610;
    wire _N10183_1612;
    wire _N10183_1613;
    wire _N10183_1615;
    wire _N10183_1622;
    wire _N10183_1623;
    wire _N10183_1624_inv;
    wire _N10183_1625;
    wire _N10183_1634;
    wire _N10183_1656;
    wire _N10183_1657;
    wire _N10183_1668;
    wire _N10183_1671;
    wire _N10183_1672;
    wire _N10183_1673;
    wire _N10183_1674;
    wire _N10183_1675;
    wire _N10183_1676;
    wire _N10183_1677;
    wire _N10183_1678;
    wire _N10183_1679;
    wire _N10183_1680;
    wire _N10183_1681;
    wire _N10183_1682;
    wire _N10183_1685;
    wire _N10183_1686;
    wire _N10183_1706;
    wire _N10183_1707;
    wire _N10183_1716;
    wire _N10183_1739;
    wire _N10183_1740;
    wire _N10183_1741;
    wire _N10183_1742;
    wire _N10183_1743;
    wire _N10183_1747;
    wire _N10183_1748;
    wire _N10183_1749;
    wire _N10183_1750;
    wire _N10183_1764;
    wire _N10183_1765;
    wire _N10183_1766;
    wire _N10183_1767;
    wire _N10183_1768;
    wire _N10183_1769;
    wire _N10183_1791;
    wire _N10183_1795;
    wire _N10183_1796;
    wire _N10183_1799;
    wire _N10183_1803;
    wire _N10183_1805;
    wire _N10183_1806;
    wire _N10183_1818;
    wire _N10183_1821;
    wire _N10183_1822;
    wire _N10183_1823;
    wire _N10183_1824;
    wire _N10183_1825;
    wire _N10183_1826;
    wire _N10183_1827;
    wire _N10183_1828;
    wire _N10183_1829;
    wire _N10183_1830;
    wire _N10183_1831;
    wire _N10183_1832;
    wire _N10183_1835;
    wire _N10183_1836;
    wire _N10183_1854;
    wire _N10183_1855;
    wire _N10183_1863;
    wire _N10183_1884;
    wire _N10183_1885;
    wire _N10183_1886;
    wire _N10183_1887;
    wire _N10183_1888;
    wire _N10183_1892;
    wire _N10183_1893;
    wire _N10183_1894;
    wire _N10183_1907;
    wire _N10183_1908;
    wire _N10183_1909;
    wire _N10183_1910;
    wire _N10183_1911;
    wire _N10183_1912;
    wire _N10183_1935;
    wire _N10183_1936;
    wire _N10183_1938;
    wire _N10183_1943;
    wire _N10183_1955;
    wire _N10183_1958;
    wire _N10183_1959;
    wire _N10183_1960;
    wire _N10183_1961;
    wire _N10183_1962;
    wire _N10183_1963;
    wire _N10183_1964;
    wire _N10183_1965;
    wire _N10183_1966;
    wire _N10183_1967;
    wire _N10183_1968;
    wire _N10183_1969;
    wire _N10183_1972;
    wire _N10183_1973;
    wire _N10183_1991;
    wire _N10183_1992;
    wire _N10183_2000;
    wire _N10183_2021;
    wire _N10183_2022;
    wire _N10183_2023;
    wire _N10183_2024;
    wire _N10183_2025;
    wire _N10183_2029;
    wire _N10183_2030;
    wire _N10183_2031;
    wire _N10183_2044;
    wire _N10183_2045;
    wire _N10183_2046;
    wire _N10183_2047;
    wire _N10183_2048;
    wire _N10183_2049;
    wire _N10183_2072;
    wire _N10183_2073;
    wire _N10183_2075;
    wire _N10183_2080;
    wire _N10183_2092;
    wire _N10183_2095;
    wire _N10183_2096;
    wire _N10183_2097;
    wire _N10183_2098;
    wire _N10183_2099;
    wire _N10183_2100;
    wire _N10183_2101;
    wire _N10183_2102;
    wire _N10183_2103;
    wire _N10183_2104;
    wire _N10183_2105;
    wire _N10183_2106;
    wire _N10183_2109;
    wire _N10183_2110;
    wire _N10183_2128;
    wire _N10183_2129;
    wire _N10183_2137;
    wire _N10183_2158;
    wire _N10183_2159;
    wire _N10183_2160;
    wire _N10183_2161;
    wire _N10183_2162;
    wire _N10183_2166;
    wire _N10183_2167;
    wire _N10183_2168;
    wire _N10183_2181;
    wire _N10183_2182;
    wire _N10183_2183;
    wire _N10183_2184;
    wire _N10183_2185;
    wire _N10183_2186;
    wire _N10183_2209;
    wire _N10183_2210;
    wire _N10183_2212;
    wire _N10183_2217;
    wire _N10183_2229;
    wire _N10183_2232;
    wire _N10183_2233;
    wire _N10183_2234;
    wire _N10183_2235;
    wire _N10183_2236;
    wire _N10183_2237;
    wire _N10183_2238;
    wire _N10183_2239;
    wire _N10183_2240;
    wire _N10183_2241;
    wire _N10183_2242;
    wire _N10183_2243;
    wire _N10183_2246;
    wire _N10183_2247;
    wire _N10183_2265;
    wire _N10183_2266;
    wire _N10183_2274;
    wire _N10183_2295;
    wire _N10183_2296;
    wire _N10183_2297;
    wire _N10183_2298;
    wire _N10183_2299;
    wire _N10183_2303;
    wire _N10183_2304;
    wire _N10183_2305;
    wire _N10183_2318;
    wire _N10183_2319;
    wire _N10183_2320;
    wire _N10183_2321;
    wire _N10183_2322;
    wire _N10183_2323;
    wire _N10183_2346;
    wire _N10183_2347;
    wire _N10183_2349;
    wire _N10183_2354;
    wire _N10183_2366;
    wire _N10183_2369;
    wire _N10183_2370;
    wire _N10183_2371;
    wire _N10183_2372;
    wire _N10183_2373;
    wire _N10183_2374;
    wire _N10183_2375;
    wire _N10183_2376;
    wire _N10183_2377;
    wire _N10183_2378;
    wire _N10183_2379;
    wire _N10183_2380;
    wire _N10183_2383;
    wire _N10183_2384;
    wire _N10183_2402;
    wire _N10183_2403;
    wire _N10183_2411;
    wire _N10183_2432;
    wire _N10183_2433;
    wire _N10183_2434;
    wire _N10183_2435;
    wire _N10183_2436;
    wire _N10183_2440;
    wire _N10183_2441;
    wire _N10183_2442;
    wire _N10183_2455;
    wire _N10183_2456;
    wire _N10183_2457;
    wire _N10183_2458;
    wire _N10183_2459;
    wire _N10183_2460;
    wire _N10183_2483;
    wire _N10183_2484;
    wire _N10183_2486;
    wire _N10183_2491;
    wire _N10183_2503;
    wire _N10183_2506;
    wire _N10183_2507;
    wire _N10183_2508;
    wire _N10183_2509;
    wire _N10183_2510;
    wire _N10183_2511;
    wire _N10183_2512;
    wire _N10183_2513;
    wire _N10183_2514;
    wire _N10183_2515;
    wire _N10183_2516;
    wire _N10183_2517;
    wire _N10183_2520;
    wire _N10183_2521;
    wire _N10183_2539;
    wire _N10183_2548;
    wire _N10183_2569;
    wire _N10183_2570;
    wire _N10183_2571;
    wire _N10183_2572;
    wire _N10183_2573;
    wire _N10183_2577;
    wire _N10183_2578;
    wire _N10183_2579;
    wire _N10183_2592;
    wire _N10183_2593;
    wire _N10183_2594;
    wire _N10183_2595;
    wire _N10183_2596;
    wire _N10183_2597;
    wire _N10183_2620;
    wire _N10183_2621;
    wire _N10183_2623;
    wire _N10183_2628;
    wire _N10183_2642;
    wire _N10183_2650;
    wire _N10183_2710;
    wire _N10183_2712;
    wire _N10183_2720;
    wire _N10183_2782;
    wire _N10183_2789;
    wire _N10183_2790;
    wire _N10183_2852;
    wire _N10183_2911;
    wire _N10183_2918;
    wire _N10183_2976;
    wire _N10183_3032;
    wire _N10183_3039;
    wire _N10183_3097;
    wire _N10183_3153;
    wire _N10183_3160;
    wire _N10183_3218;
    wire _N10183_3274;
    wire _N10183_3281;
    wire _N10183_3339;
    wire _N10183_3395;
    wire _N10183_3402;
    wire _N10183_3460;
    wire _N10183_3516;
    wire _N10183_3523;
    wire _N10183_3556;
    wire _N10233;
    wire _N10246;
    wire _N10315;
    wire _N10344;
    wire _N10345;
    wire _N10361;
    wire _N10441;
    wire _N10456;
    wire _N10457;
    wire _N10481;
    wire _N10483;
    wire _N10495;
    wire _N10496;
    wire _N10499;
    wire _N10500;
    wire _N10501;
    wire _N10502;
    wire _N10505;
    wire _N10511;
    wire _N10517;
    wire _N10518;
    wire _N10519;
    wire _N10520;
    wire _N10521;
    wire _N10526;
    wire _N10532;
    wire _N10539;
    wire _N10540;
    wire _N10545;
    wire _N10546;
    wire _N10547;
    wire _N10548;
    wire _N10558;
    wire _N10560;
    wire _N10566;
    wire _N10567;
    wire _N10568;
    wire _N10569;
    wire _N10570;
    wire _N10571;
    wire _N10580;
    wire _N10584;
    wire _N10585;
    wire _N10592;
    wire _N10844;
    wire _N10904_2;
    wire _N10911_2;
    wire _N10911_3;
    wire _N10924_2;
    wire _N10992_1;
    wire _N10992_3;
    wire _N11004_2;
    wire _N11014_3;
    wire _N11016_2;
    wire _N11036_2;
    wire _N11036_3;
    wire _N11162_2;
    wire _N11162_3;
    wire _N11168_2;
    wire _N11179_2;
    wire _N11190_2;
    wire _N11198_2;
    wire _N11198_5;
    wire _N11198_6;
    wire _N11227_2;
    wire _N11227_3;
    wire _N11259_2;
    wire _N11259_3;
    wire _N11319_2;
    wire _N11364_2;
    wire _N11426_3;
    wire _N11428_2;
    wire _N11428_3;
    wire _N11482_2;
    wire _N11482_3;
    wire _N11489_2;
    wire _N11502_2;
    wire _N11503_2;
    wire _N11792_3;
    wire _N11805;
    wire _N11806;
    wire _N11807;
    wire _N11808;
    wire _N11809;
    wire _N11810;
    wire _N11811;
    wire _N11812;
    wire _N11813;
    wire _N11814;
    wire _N11824;
    wire _N11834;
    wire _N11839;
    wire _N11860;
    wire _N11868;
    wire _N11882;
    wire _N11890;
    wire _N11897;
    wire _N11899;
    wire _N11901;
    wire _N11905;
    wire _N11914;
    wire _N11923;
    wire _N11925;
    wire _N11928;
    wire _N11935;
    wire _N11940;
    wire _N11945;
    wire _N11956;
    wire _N11958;
    wire _N11960;
    wire _N11966;
    wire _N11968;
    wire _N11972;
    wire _N11979;
    wire _N11987;
    wire _N11990;
    wire _N11998;
    wire _N12002;
    wire _N12010;
    wire _N12012;
    wire _N12013;
    wire _N12029;
    wire _N12037;
    wire _N12039;
    wire _N12050;
    wire _N12065;
    wire _N12187;
    wire _N12189;
    wire _N12192;
    wire _N12199;
    wire _N12216;
    wire _N12219;
    wire _N12220;
    wire _N12225;
    wire _N12226;
    wire _N12227;
    wire _N12228;
    wire _N12229;
    wire _N12230;
    wire _N12231;
    wire _N12282;
    wire _N12284;
    wire _N12286;
    wire _N12288;
    wire _N12290;
    wire _N12292;
    wire _N12294;
    wire _N12317;
    wire [31:0] data;
    wire [15:0] lcd_id;
    wire nt_lcd_clk;
    wire nt_lcd_de;
    wire nt_lcd_de_inv;
    wire nt_sys_clk;
    wire nt_sys_rst_n;
    wire nt_touch_rst_n;
    wire nt_touch_scl;
    wire [15:0] \u_lcd_rgb_char/bcd_data_x ;
    wire [15:0] \u_lcd_rgb_char/bcd_data_y ;
    wire [23:0] \u_lcd_rgb_char/lcd_rgb_o ;
    wire [23:0] \u_lcd_rgb_char/pixel_data_w ;
    wire [10:0] \u_lcd_rgb_char/pixel_xpos_w ;
    wire [10:0] \u_lcd_rgb_char/pixel_ypos_w ;
    wire \u_lcd_rgb_char/pixel_ypos_w[0]_inv ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N0 ;
    wire [4:0] \u_lcd_rgb_char/u_binary2bcd_x/N7 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N19 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N23 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N31 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N39 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N47 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N73 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N76 ;
    wire [4:0] \u_lcd_rgb_char/u_binary2bcd_x/N90 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N94 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N95 ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/N97 ;
    wire [3:0] \u_lcd_rgb_char/u_binary2bcd_x/N98 ;
    wire [3:0] \u_lcd_rgb_char/u_binary2bcd_x/N104 ;
    wire [3:0] \u_lcd_rgb_char/u_binary2bcd_x/N110 ;
    wire [3:0] \u_lcd_rgb_char/u_binary2bcd_x/N116 ;
    wire [14:0] \u_lcd_rgb_char/u_binary2bcd_x/N122 ;
    wire [4:0] \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift ;
    wire [31:0] \u_lcd_rgb_char/u_binary2bcd_x/data_shift ;
    wire \u_lcd_rgb_char/u_binary2bcd_x/shift_flag ;
    wire [4:0] \u_lcd_rgb_char/u_binary2bcd_y/N7 ;
    wire \u_lcd_rgb_char/u_binary2bcd_y/N23 ;
    wire \u_lcd_rgb_char/u_binary2bcd_y/N31 ;
    wire \u_lcd_rgb_char/u_binary2bcd_y/N39 ;
    wire \u_lcd_rgb_char/u_binary2bcd_y/N73 ;
    wire \u_lcd_rgb_char/u_binary2bcd_y/N76 ;
    wire [4:0] \u_lcd_rgb_char/u_binary2bcd_y/N90 ;
    wire \u_lcd_rgb_char/u_binary2bcd_y/N94 ;
    wire \u_lcd_rgb_char/u_binary2bcd_y/N95 ;
    wire \u_lcd_rgb_char/u_binary2bcd_y/N97 ;
    wire [3:0] \u_lcd_rgb_char/u_binary2bcd_y/N104 ;
    wire [3:0] \u_lcd_rgb_char/u_binary2bcd_y/N110 ;
    wire [3:0] \u_lcd_rgb_char/u_binary2bcd_y/N116 ;
    wire [14:0] \u_lcd_rgb_char/u_binary2bcd_y/N122 ;
    wire [4:0] \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift ;
    wire [31:0] \u_lcd_rgb_char/u_binary2bcd_y/data_shift ;
    wire \u_lcd_rgb_char/u_clk_div/N3 ;
    wire \u_lcd_rgb_char/u_clk_div/N39 ;
    wire \u_lcd_rgb_char/u_clk_div/N40 ;
    wire \u_lcd_rgb_char/u_clk_div/clk_12_5m ;
    wire \u_lcd_rgb_char/u_clk_div/div_4_cnt ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_display/N46_1.co ;
    wire [31:0] \u_lcd_rgb_char/u_lcd_display/N59 ;
    wire [13:0] \u_lcd_rgb_char/u_lcd_display/N59_1.co ;
    wire [35:0] \u_lcd_rgb_char/u_lcd_display/N392 ;
    wire [23:0] \u_lcd_rgb_char/u_lcd_display/N9971 ;
    wire [11:0] \u_lcd_rgb_char/u_lcd_driver/N7_1.co ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N7_4.co ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N12 ;
    wire \u_lcd_rgb_char/u_lcd_driver/N13 ;
    wire [11:0] \u_lcd_rgb_char/u_lcd_driver/N13.co ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N16 ;
    wire \u_lcd_rgb_char/u_lcd_driver/N17 ;
    wire [11:0] \u_lcd_rgb_char/u_lcd_driver/N17.co ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N23 ;
    wire [11:0] \u_lcd_rgb_char/u_lcd_driver/N25.co ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N98 ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N100 ;
    wire [8:0] \u_lcd_rgb_char/u_lcd_driver/N100_1.co ;
    wire \u_lcd_rgb_char/u_lcd_driver/N101 ;
    wire [11:0] \u_lcd_rgb_char/u_lcd_driver/N101.co ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N106 ;
    wire \u_lcd_rgb_char/u_lcd_driver/N107 ;
    wire [11:0] \u_lcd_rgb_char/u_lcd_driver/N107.co ;
    wire \u_lcd_rgb_char/u_lcd_driver/N116 ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N124 ;
    wire [6:0] \u_lcd_rgb_char/u_lcd_driver/N124_1.co ;
    wire \u_lcd_rgb_char/u_lcd_driver/N125 ;
    wire [11:0] \u_lcd_rgb_char/u_lcd_driver/N125.co ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N144 ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N144_1.co ;
    wire \u_lcd_rgb_char/u_lcd_driver/N145 ;
    wire [11:0] \u_lcd_rgb_char/u_lcd_driver/N145.co ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N153 ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N178 ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N180 ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/N182 ;
    wire \u_lcd_rgb_char/u_lcd_driver/data_req ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/h_back ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/h_cnt ;
    wire \u_lcd_rgb_char/u_lcd_driver/h_cnt[1]_inv ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/h_disp ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/h_sync ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/h_total ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/nb0 ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/nb1 ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/nb3 ;
    wire [10:0] \u_lcd_rgb_char/u_lcd_driver/v_cnt ;
    wire \u_lcd_rgb_char/u_lcd_driver/v_cnt[0]_inv ;
    wire [15:0] \u_lcd_rgb_char/u_rd_id/N22 ;
    wire \u_lcd_rgb_char/u_rd_id/N27 ;
    wire \u_lcd_rgb_char/u_rd_id/N31 ;
    wire \u_lcd_rgb_char/u_rd_id/N35 ;
    wire \u_lcd_rgb_char/u_rd_id/rd_flag ;
    wire \u_touch_top/bit_ctrl ;
    wire \u_touch_top/dri_clk ;
    wire \u_touch_top/i2c_ack ;
    wire [15:0] \u_touch_top/i2c_addr ;
    wire [7:0] \u_touch_top/i2c_data_r ;
    wire [7:0] \u_touch_top/i2c_data_w ;
    wire \u_touch_top/i2c_done ;
    wire \u_touch_top/i2c_exec ;
    wire \u_touch_top/i2c_rh_wl ;
    wire \u_touch_top/once_byte_done ;
    wire [7:0] \u_touch_top/reg_num ;
    wire [6:0] \u_touch_top/slave_addr ;
    wire [8:0] \u_touch_top/u_i2c_dri/N2.co ;
    wire [9:0] \u_touch_top/u_i2c_dri/N12 ;
    wire [6:0] \u_touch_top/u_i2c_dri/N97 ;
    wire [7:0] \u_touch_top/u_i2c_dri/N475 ;
    wire [7:0] \u_touch_top/u_i2c_dri/N475_1.co ;
    wire \u_touch_top/u_i2c_dri/N476 ;
    wire [8:0] \u_touch_top/u_i2c_dri/N476.co ;
    wire [6:0] \u_touch_top/u_i2c_dri/N552 ;
    wire \u_touch_top/u_i2c_dri/N557 ;
    wire \u_touch_top/u_i2c_dri/N558 ;
    wire \u_touch_top/u_i2c_dri/N582_inv ;
    wire \u_touch_top/u_i2c_dri/N607 ;
    wire \u_touch_top/u_i2c_dri/N637 ;
    wire [9:0] \u_touch_top/u_i2c_dri/N811 ;
    wire \u_touch_top/u_i2c_dri/N814 ;
    wire [7:0] \u_touch_top/u_i2c_dri/N815 ;
    wire \u_touch_top/u_i2c_dri/N1180 ;
    wire \u_touch_top/u_i2c_dri/N1185 ;
    wire \u_touch_top/u_i2c_dri/N1222 ;
    wire \u_touch_top/u_i2c_dri/N1227 ;
    wire \u_touch_top/u_i2c_dri/N1230 ;
    wire \u_touch_top/u_i2c_dri/N1232 ;
    wire \u_touch_top/u_i2c_dri/N1600 ;
    wire \u_touch_top/u_i2c_dri/N1668 ;
    wire \u_touch_top/u_i2c_dri/N2082 ;
    wire \u_touch_top/u_i2c_dri/N2434 ;
    wire \u_touch_top/u_i2c_dri/N2868 ;
    wire \u_touch_top/u_i2c_dri/N2917 ;
    wire \u_touch_top/u_i2c_dri/N2925 ;
    wire \u_touch_top/u_i2c_dri/N3005 ;
    wire \u_touch_top/u_i2c_dri/N3052 ;
    wire \u_touch_top/u_i2c_dri/N3102 ;
    wire \u_touch_top/u_i2c_dri/N3152 ;
    wire \u_touch_top/u_i2c_dri/N3202 ;
    wire \u_touch_top/u_i2c_dri/N3252 ;
    wire \u_touch_top/u_i2c_dri/N3302 ;
    wire \u_touch_top/u_i2c_dri/N3352 ;
    wire \u_touch_top/u_i2c_dri/_N2 ;
    wire \u_touch_top/u_i2c_dri/_N5 ;
    wire \u_touch_top/u_i2c_dri/_N9 ;
    wire \u_touch_top/u_i2c_dri/_N15 ;
    wire \u_touch_top/u_i2c_dri/_N19 ;
    wire \u_touch_top/u_i2c_dri/_N23 ;
    wire \u_touch_top/u_i2c_dri/_N27 ;
    wire \u_touch_top/u_i2c_dri/_N39 ;
    wire \u_touch_top/u_i2c_dri/_N42 ;
    wire [15:0] \u_touch_top/u_i2c_dri/addr_t ;
    wire [9:0] \u_touch_top/u_i2c_dri/clk_cnt ;
    wire \u_touch_top/u_i2c_dri/clk_cnt[0]_inv ;
    wire [6:0] \u_touch_top/u_i2c_dri/cnt ;
    wire [7:0] \u_touch_top/u_i2c_dri/cur_state_reg ;
    wire [7:0] \u_touch_top/u_i2c_dri/data_r ;
    wire [7:0] \u_touch_top/u_i2c_dri/data_wr_t ;
    wire [7:0] \u_touch_top/u_i2c_dri/reg_cnt ;
    wire \u_touch_top/u_i2c_dri/reg_done ;
    wire \u_touch_top/u_i2c_dri/sda_dir ;
    wire \u_touch_top/u_i2c_dri/sda_dir_inv ;
    wire \u_touch_top/u_i2c_dri/sda_out ;
    wire \u_touch_top/u_i2c_dri/st_done ;
    wire \u_touch_top/u_i2c_dri/wr_flag ;
    wire \u_touch_top/u_touch_dri/N70 ;
    wire \u_touch_top/u_touch_dri/N166 ;
    wire \u_touch_top/u_touch_dri/N296 ;
    wire [15:0] \u_touch_top/u_touch_dri/N376 ;
    wire [15:0] \u_touch_top/u_touch_dri/N377 ;
    wire \u_touch_top/u_touch_dri/N390 ;
    wire \u_touch_top/u_touch_dri/N394 ;
    wire \u_touch_top/u_touch_dri/N474 ;
    wire [19:0] \u_touch_top/u_touch_dri/N559 ;
    wire \u_touch_top/u_touch_dri/N614 ;
    wire \u_touch_top/u_touch_dri/N641 ;
    wire \u_touch_top/u_touch_dri/N642 ;
    wire \u_touch_top/u_touch_dri/N666 ;
    wire \u_touch_top/u_touch_dri/N716 ;
    wire \u_touch_top/u_touch_dri/N739 ;
    wire \u_touch_top/u_touch_dri/N863 ;
    wire \u_touch_top/u_touch_dri/N905 ;
    wire \u_touch_top/u_touch_dri/N924 ;
    wire \u_touch_top/u_touch_dri/N933 ;
    wire \u_touch_top/u_touch_dri/N935 ;
    wire \u_touch_top/u_touch_dri/N937 ;
    wire \u_touch_top/u_touch_dri/N944 ;
    wire \u_touch_top/u_touch_dri/N945 ;
    wire \u_touch_top/u_touch_dri/N948 ;
    wire \u_touch_top/u_touch_dri/N961 ;
    wire \u_touch_top/u_touch_dri/N1074 ;
    wire \u_touch_top/u_touch_dri/N1201 ;
    wire \u_touch_top/u_touch_dri/N1206 ;
    wire \u_touch_top/u_touch_dri/N1216 ;
    wire \u_touch_top/u_touch_dri/N1218 ;
    wire \u_touch_top/u_touch_dri/N1281 ;
    wire \u_touch_top/u_touch_dri/N1297 ;
    wire [15:0] \u_touch_top/u_touch_dri/N1300 ;
    wire \u_touch_top/u_touch_dri/N1450 ;
    wire \u_touch_top/u_touch_dri/N1453 ;
    wire \u_touch_top/u_touch_dri/N1494 ;
    wire \u_touch_top/u_touch_dri/N1497 ;
    wire \u_touch_top/u_touch_dri/N1529 ;
    wire \u_touch_top/u_touch_dri/N1569 ;
    wire \u_touch_top/u_touch_dri/N1610 ;
    wire [9:0] \u_touch_top/u_touch_dri/N1629 ;
    wire \u_touch_top/u_touch_dri/_N48 ;
    wire \u_touch_top/u_touch_dri/_N51 ;
    wire \u_touch_top/u_touch_dri/_N55 ;
    wire \u_touch_top/u_touch_dri/_N61 ;
    wire \u_touch_top/u_touch_dri/_N64 ;
    wire \u_touch_top/u_touch_dri/_N67 ;
    wire \u_touch_top/u_touch_dri/_N70 ;
    wire \u_touch_top/u_touch_dri/_N74 ;
    wire \u_touch_top/u_touch_dri/_N81 ;
    wire \u_touch_top/u_touch_dri/_N85 ;
    wire \u_touch_top/u_touch_dri/_N91 ;
    wire \u_touch_top/u_touch_dri/_N95 ;
    wire \u_touch_top/u_touch_dri/_N99 ;
    wire \u_touch_top/u_touch_dri/_N102 ;
    wire \u_touch_top/u_touch_dri/_N107 ;
    wire \u_touch_top/u_touch_dri/_N111 ;
    wire \u_touch_top/u_touch_dri/_N119 ;
    wire \u_touch_top/u_touch_dri/_N120 ;
    wire \u_touch_top/u_touch_dri/_N126 ;
    wire \u_touch_top/u_touch_dri/_N131 ;
    wire [15:0] \u_touch_top/u_touch_dri/chip_version ;
    wire [19:0] \u_touch_top/u_touch_dri/cnt_time ;
    wire \u_touch_top/u_touch_dri/cnt_time_en ;
    wire [15:0] \u_touch_top/u_touch_dri/coord_reg ;
    wire [6:0] \u_touch_top/u_touch_dri/cur_state_reg ;
    wire [7:0] \u_touch_top/u_touch_dri/flow_cnt_reg ;
    wire \u_touch_top/u_touch_dri/ft_flag ;
    wire [6:0] \u_touch_top/u_touch_dri/next_state ;
    wire \u_touch_top/u_touch_dri/st_done ;
    wire \u_touch_top/u_touch_dri/touch_int_dir ;
    wire \u_touch_top/u_touch_dri/touch_int_dir_inv ;
    wire \u_touch_top/u_touch_dri/touch_int_out ;
    wire [15:0] \u_touch_top/u_touch_dri/touch_s_reg ;
    wire \u_touch_top/u_touch_dri/touch_valid ;
    wire [15:0] \u_touch_top/u_touch_dri/tp_x_coord ;
    wire [15:0] \u_touch_top/u_touch_dri/tp_x_coord_t ;
    wire [15:0] \u_touch_top/u_touch_dri/tp_y_coord ;
    wire [15:0] \u_touch_top/u_touch_dri/tp_y_coord_t ;

    GTP_GRS GRS_INST (
            .GRS_N (1'b1));

    GTP_LUT5M /* _N10183_87_inv */ #(
            .INIT(32'b00010001110111011110001011100010))
        _N10183_87_inv_vname (
            .Z (_N10183_87_inv),
            .I0 (_N10183_250),
            .I1 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I2 (_N10183_251),
            .I3 (_N10183_252),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (_N10183_249));
    // defparam _N10183_87_inv_vname.orig_name = _N10183_87_inv;
	// LUT = (I1&I2&~I4)|(ID&~I1&~I4)|(I1&~I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5M /* _N10183_91_inv */ #(
            .INIT(32'b00010001110111011110001011100010))
        _N10183_91_inv_vname (
            .Z (_N10183_91_inv),
            .I0 (_N10183_266),
            .I1 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I2 (_N10183_267),
            .I3 (_N10183_268),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (_N10183_265));
    // defparam _N10183_91_inv_vname.orig_name = _N10183_91_inv;
	// LUT = (I1&I2&~I4)|(ID&~I1&~I4)|(I1&~I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5M /* _N10183_95_inv */ #(
            .INIT(32'b00010001110111011110001011100010))
        _N10183_95_inv_vname (
            .Z (_N10183_95_inv),
            .I0 (_N10183_282),
            .I1 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I2 (_N10183_283),
            .I3 (_N10183_284),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (_N10183_281));
    // defparam _N10183_95_inv_vname.orig_name = _N10183_95_inv;
	// LUT = (I1&I2&~I4)|(ID&~I1&~I4)|(I1&~I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5M /* _N10183_319_inv */ #(
            .INIT(32'b00011011000110111111101000001010))
        _N10183_319_inv_vname (
            .Z (_N10183_319_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (_N10183_1028),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (_N10183_1030),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (_N10183_1029));
    // defparam _N10183_319_inv_vname.orig_name = _N10183_319_inv;
	// LUT = (I2&I3&~I4)|(ID&~I2&~I4)|(I0&~I2&I4)|(~I0&~I1&I4) ;

    GTP_LUT4 /* _N10183_323_inv */ #(
            .INIT(16'b0111001011111010))
        _N10183_323_inv_vname (
            .Z (_N10183_323_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (_N10183_589),
            .I3 (_N10183_1043));
    // defparam _N10183_323_inv_vname.orig_name = _N10183_323_inv;
	// LUT = (I0&~I3)|(~I0&I2)|(I0&~I1) ;

    GTP_LUT5M /* _N10183_331_inv */ #(
            .INIT(32'b01010001000100011010101010101010))
        _N10183_331_inv_vname (
            .Z (_N10183_331_inv),
            .I0 (_N10183_1064),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_2720),
            .I4 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .ID (_N10183_602));
    // defparam _N10183_331_inv_vname.orig_name = _N10183_331_inv;
	// LUT = (ID&~I4)|(~I0&I2&I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5M /* _N10183_350_inv */ #(
            .INIT(32'b00011011000110111111101000001010))
        _N10183_350_inv_vname (
            .Z (_N10183_350_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (_N10183_1121),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (_N10183_1123),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (_N10183_1122));
    // defparam _N10183_350_inv_vname.orig_name = _N10183_350_inv;
	// LUT = (I2&I3&~I4)|(ID&~I2&~I4)|(I0&~I2&I4)|(~I0&~I1&I4) ;

    GTP_LUT4 /* _N10183_354_inv */ #(
            .INIT(16'b0111001011111010))
        _N10183_354_inv_vname (
            .Z (_N10183_354_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (_N10183_645),
            .I3 (_N10183_1136));
    // defparam _N10183_354_inv_vname.orig_name = _N10183_354_inv;
	// LUT = (I0&~I3)|(~I0&I2)|(I0&~I1) ;

    GTP_LUT5M /* _N10183_362_inv */ #(
            .INIT(32'b01010001000100011010101010101010))
        _N10183_362_inv_vname (
            .Z (_N10183_362_inv),
            .I0 (_N10183_1064),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_2720),
            .I4 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .ID (_N10183_658));
    // defparam _N10183_362_inv_vname.orig_name = _N10183_362_inv;
	// LUT = (ID&~I4)|(~I0&I2&I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5M /* _N10183_381_inv */ #(
            .INIT(32'b00011011000110111111101000001010))
        _N10183_381_inv_vname (
            .Z (_N10183_381_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (_N10183_1212),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (_N10183_1214),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (_N10183_1213));
    // defparam _N10183_381_inv_vname.orig_name = _N10183_381_inv;
	// LUT = (I2&I3&~I4)|(ID&~I2&~I4)|(I0&~I2&I4)|(~I0&~I1&I4) ;

    GTP_LUT4 /* _N10183_385_inv */ #(
            .INIT(16'b0111001011111010))
        _N10183_385_inv_vname (
            .Z (_N10183_385_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (_N10183_701),
            .I3 (_N10183_1227));
    // defparam _N10183_385_inv_vname.orig_name = _N10183_385_inv;
	// LUT = (I0&~I3)|(~I0&I2)|(I0&~I1) ;

    GTP_LUT5M /* _N10183_393_inv */ #(
            .INIT(32'b01010001000100011010101010101010))
        _N10183_393_inv_vname (
            .Z (_N10183_393_inv),
            .I0 (_N10183_1064),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_2720),
            .I4 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .ID (_N10183_714));
    // defparam _N10183_393_inv_vname.orig_name = _N10183_393_inv;
	// LUT = (ID&~I4)|(~I0&I2&I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5M /* _N10183_412_inv */ #(
            .INIT(32'b00011011000110111111101000001010))
        _N10183_412_inv_vname (
            .Z (_N10183_412_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (_N10183_1303),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (_N10183_1305),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (_N10183_1304));
    // defparam _N10183_412_inv_vname.orig_name = _N10183_412_inv;
	// LUT = (I2&I3&~I4)|(ID&~I2&~I4)|(I0&~I2&I4)|(~I0&~I1&I4) ;

    GTP_LUT4 /* _N10183_416_inv */ #(
            .INIT(16'b0111001011111010))
        _N10183_416_inv_vname (
            .Z (_N10183_416_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (_N10183_757),
            .I3 (_N10183_1318));
    // defparam _N10183_416_inv_vname.orig_name = _N10183_416_inv;
	// LUT = (I0&~I3)|(~I0&I2)|(I0&~I1) ;

    GTP_LUT5M /* _N10183_424_inv */ #(
            .INIT(32'b01010001000100011010101010101010))
        _N10183_424_inv_vname (
            .Z (_N10183_424_inv),
            .I0 (_N10183_1064),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_2720),
            .I4 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .ID (_N10183_770));
    // defparam _N10183_424_inv_vname.orig_name = _N10183_424_inv;
	// LUT = (ID&~I4)|(~I0&I2&I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5M /* _N10183_443_inv */ #(
            .INIT(32'b00011011000110111111101000001010))
        _N10183_443_inv_vname (
            .Z (_N10183_443_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (_N10183_1394),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (_N10183_1396),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (_N10183_1395));
    // defparam _N10183_443_inv_vname.orig_name = _N10183_443_inv;
	// LUT = (I2&I3&~I4)|(ID&~I2&~I4)|(I0&~I2&I4)|(~I0&~I1&I4) ;

    GTP_LUT4 /* _N10183_447_inv */ #(
            .INIT(16'b0111001011111010))
        _N10183_447_inv_vname (
            .Z (_N10183_447_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (_N10183_813),
            .I3 (_N10183_1409));
    // defparam _N10183_447_inv_vname.orig_name = _N10183_447_inv;
	// LUT = (I0&~I3)|(~I0&I2)|(I0&~I1) ;

    GTP_LUT5M /* _N10183_455_inv */ #(
            .INIT(32'b01010001000100011010101010101010))
        _N10183_455_inv_vname (
            .Z (_N10183_455_inv),
            .I0 (_N10183_1064),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_2720),
            .I4 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .ID (_N10183_826));
    // defparam _N10183_455_inv_vname.orig_name = _N10183_455_inv;
	// LUT = (ID&~I4)|(~I0&I2&I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5M /* _N10183_474_inv */ #(
            .INIT(32'b00011011000110111111101000001010))
        _N10183_474_inv_vname (
            .Z (_N10183_474_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (_N10183_1485),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (_N10183_1487),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (_N10183_1486));
    // defparam _N10183_474_inv_vname.orig_name = _N10183_474_inv;
	// LUT = (I2&I3&~I4)|(ID&~I2&~I4)|(I0&~I2&I4)|(~I0&~I1&I4) ;

    GTP_LUT4 /* _N10183_478_inv */ #(
            .INIT(16'b0111001011111010))
        _N10183_478_inv_vname (
            .Z (_N10183_478_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (_N10183_869),
            .I3 (_N10183_1500));
    // defparam _N10183_478_inv_vname.orig_name = _N10183_478_inv;
	// LUT = (I0&~I3)|(~I0&I2)|(I0&~I1) ;

    GTP_LUT5M /* _N10183_486_inv */ #(
            .INIT(32'b01010001000100011010101010101010))
        _N10183_486_inv_vname (
            .Z (_N10183_486_inv),
            .I0 (_N10183_1064),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_2720),
            .I4 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .ID (_N10183_882));
    // defparam _N10183_486_inv_vname.orig_name = _N10183_486_inv;
	// LUT = (ID&~I4)|(~I0&I2&I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5M /* _N10183_505_inv */ #(
            .INIT(32'b00011011000110111111101000001010))
        _N10183_505_inv_vname (
            .Z (_N10183_505_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (_N10183_1576),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (_N10183_1578),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (_N10183_1577));
    // defparam _N10183_505_inv_vname.orig_name = _N10183_505_inv;
	// LUT = (I2&I3&~I4)|(ID&~I2&~I4)|(I0&~I2&I4)|(~I0&~I1&I4) ;

    GTP_LUT4 /* _N10183_509_inv */ #(
            .INIT(16'b0111001011111010))
        _N10183_509_inv_vname (
            .Z (_N10183_509_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (_N10183_925),
            .I3 (_N10183_1591));
    // defparam _N10183_509_inv_vname.orig_name = _N10183_509_inv;
	// LUT = (I0&~I3)|(~I0&I2)|(I0&~I1) ;

    GTP_LUT5M /* _N10183_517_inv */ #(
            .INIT(32'b01010001000100011010101010101010))
        _N10183_517_inv_vname (
            .Z (_N10183_517_inv),
            .I0 (_N10183_1064),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_2720),
            .I4 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .ID (_N10183_938));
    // defparam _N10183_517_inv_vname.orig_name = _N10183_517_inv;
	// LUT = (ID&~I4)|(~I0&I2&I3&I4)|(~I0&~I1&I4) ;

    GTP_LUT5 /* _N10183_574_inv */ #(
            .INIT(32'b00100010111111010110011011111101))
        _N10183_574_inv_vname (
            .Z (_N10183_574_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_2712));
    // defparam _N10183_574_inv_vname.orig_name = _N10183_574_inv;
	// LUT = (~I0&I1&~I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_631_inv */ #(
            .INIT(32'b00100010111111010110011011111101))
        _N10183_631_inv_vname (
            .Z (_N10183_631_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_2712));
    // defparam _N10183_631_inv_vname.orig_name = _N10183_631_inv;
	// LUT = (~I0&I1&~I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_687_inv */ #(
            .INIT(32'b00100010111111010110011011111101))
        _N10183_687_inv_vname (
            .Z (_N10183_687_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_2712));
    // defparam _N10183_687_inv_vname.orig_name = _N10183_687_inv;
	// LUT = (~I0&I1&~I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_743_inv */ #(
            .INIT(32'b00100010111111010110011011111101))
        _N10183_743_inv_vname (
            .Z (_N10183_743_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_2712));
    // defparam _N10183_743_inv_vname.orig_name = _N10183_743_inv;
	// LUT = (~I0&I1&~I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_799_inv */ #(
            .INIT(32'b00100010111111010110011011111101))
        _N10183_799_inv_vname (
            .Z (_N10183_799_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_2712));
    // defparam _N10183_799_inv_vname.orig_name = _N10183_799_inv;
	// LUT = (~I0&I1&~I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_855_inv */ #(
            .INIT(32'b00100010111111010110011011111101))
        _N10183_855_inv_vname (
            .Z (_N10183_855_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_2712));
    // defparam _N10183_855_inv_vname.orig_name = _N10183_855_inv;
	// LUT = (~I0&I1&~I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_911_inv */ #(
            .INIT(32'b00100010111111010110011011111101))
        _N10183_911_inv_vname (
            .Z (_N10183_911_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_2712));
    // defparam _N10183_911_inv_vname.orig_name = _N10183_911_inv;
	// LUT = (~I0&I1&~I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_985_inv */ #(
            .INIT(32'b00000101001001000010010011011111))
        _N10183_985_inv_vname (
            .Z (_N10183_985_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
    // defparam _N10183_985_inv_vname.orig_name = _N10183_985_inv;
	// LUT = (~I2&~I3&~I4)|(I1&~I3&~I4)|(~I0&~I3&~I4)|(I0&~I1&I2&I3&~I4)|(I0&~I1&I2&~I3&I4)|(~I0&~I2&I3&I4)|(~I0&I1&~I2) ;

    GTP_LUT5 /* _N10183_1001_inv */ #(
            .INIT(32'b00011100110100100100000011100110))
        _N10183_1001_inv_vname (
            .Z (_N10183_1001_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1001_inv_vname.orig_name = _N10183_1001_inv;
	// LUT = (I0&~I1&~I3&~I4)|(~I0&I1&~I3&~I4)|(~I0&I1&I2&~I4)|(I1&~I2&I3&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(I1&I2&~I3) ;

    GTP_LUT5 /* _N10183_1011_inv */ #(
            .INIT(32'b01111111011111110011011110110111))
        _N10183_1011_inv_vname (
            .Z (_N10183_1011_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1011_inv_vname.orig_name = _N10183_1011_inv;
	// LUT = (I0&I2&~I3&~I4)|(~I2&I4)|(~I0&I4)|(~I0&~I2)|(~I1) ;

    GTP_LUT5 /* _N10183_1020_inv */ #(
            .INIT(32'b01100110111111010011011011111101))
        _N10183_1020_inv_vname (
            .Z (_N10183_1020_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1020_inv_vname.orig_name = _N10183_1020_inv;
	// LUT = (~I1&I2&~I4)|(~I0&I1&I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(~I0&I1&~I2)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_1022_inv */ #(
            .INIT(32'b00000000110111110000000000000010))
        _N10183_1022_inv_vname (
            .Z (_N10183_1022_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1022_inv_vname.orig_name = _N10183_1022_inv;
	// LUT = (I1&~I3&I4)|(~I0&~I3&I4)|(I0&~I1&~I2&~I3) ;

    GTP_LUT5 /* _N10183_1058_inv */ #(
            .INIT(32'b01010111010001111100111111100111))
        _N10183_1058_inv_vname (
            .Z (_N10183_1058_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1058_inv_vname.orig_name = _N10183_1058_inv;
	// LUT = (I0&~I1&~I3&~I4)|(I1&I3&~I4)|(I1&I2&~I4)|(~I0&I3&I4)|(~I1&~I2)|(~I0&I1) ;

    GTP_LUT5M /* _N10183_1062_inv */ #(
            .INIT(32'b00000000000000100011111011001100))
        _N10183_1062_inv_vname (
            .Z (_N10183_1062_inv),
            .I0 (_N10183_3556),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1062_inv_vname.orig_name = _N10183_1062_inv;
	// LUT = (I1&~I3&~I4)|(~I1&I2&I3&~I4)|(ID&~I1&I3&~I4)|(I1&~I2&~I4)|(I0&~I1&~I2&~I3&I4) ;

    GTP_LUT5 /* _N10183_1078_inv */ #(
            .INIT(32'b00010111011101111111000111111111))
        _N10183_1078_inv_vname (
            .Z (_N10183_1078_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1078_inv_vname.orig_name = _N10183_1078_inv;
	// LUT = (~I3&~I4)|(I2&~I4)|(~I1&~I2&I4)|(~I0&~I2&I4)|(~I1&~I3)|(~I0&~I3)|(~I0&~I1) ;

    GTP_LUT5 /* _N10183_1081_inv */ #(
            .INIT(32'b00000101001001000010010011011111))
        _N10183_1081_inv_vname (
            .Z (_N10183_1081_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
    // defparam _N10183_1081_inv_vname.orig_name = _N10183_1081_inv;
	// LUT = (~I2&~I3&~I4)|(I1&~I3&~I4)|(~I0&~I3&~I4)|(I0&~I1&I2&I3&~I4)|(I0&~I1&I2&~I3&I4)|(~I0&~I2&I3&I4)|(~I0&I1&~I2) ;

    GTP_LUT5 /* _N10183_1097_inv */ #(
            .INIT(32'b00011100110100100100000011100110))
        _N10183_1097_inv_vname (
            .Z (_N10183_1097_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1097_inv_vname.orig_name = _N10183_1097_inv;
	// LUT = (I0&~I1&~I3&~I4)|(~I0&I1&~I3&~I4)|(~I0&I1&I2&~I4)|(I1&~I2&I3&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(I1&I2&~I3) ;

    GTP_LUT5 /* _N10183_1104_inv */ #(
            .INIT(32'b01111111011111110011011110110111))
        _N10183_1104_inv_vname (
            .Z (_N10183_1104_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1104_inv_vname.orig_name = _N10183_1104_inv;
	// LUT = (I0&I2&~I3&~I4)|(~I2&I4)|(~I0&I4)|(~I0&~I2)|(~I1) ;

    GTP_LUT5 /* _N10183_1113_inv */ #(
            .INIT(32'b01100110111111010011011011111101))
        _N10183_1113_inv_vname (
            .Z (_N10183_1113_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1113_inv_vname.orig_name = _N10183_1113_inv;
	// LUT = (~I1&I2&~I4)|(~I0&I1&I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(~I0&I1&~I2)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_1115_inv */ #(
            .INIT(32'b00000000110111110000000000000010))
        _N10183_1115_inv_vname (
            .Z (_N10183_1115_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1115_inv_vname.orig_name = _N10183_1115_inv;
	// LUT = (I1&~I3&I4)|(~I0&~I3&I4)|(I0&~I1&~I2&~I3) ;

    GTP_LUT5 /* _N10183_1150_inv */ #(
            .INIT(32'b01010111010001111100111111100111))
        _N10183_1150_inv_vname (
            .Z (_N10183_1150_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1150_inv_vname.orig_name = _N10183_1150_inv;
	// LUT = (I0&~I1&~I3&~I4)|(I1&I3&~I4)|(I1&I2&~I4)|(~I0&I3&I4)|(~I1&~I2)|(~I0&I1) ;

    GTP_LUT5M /* _N10183_1154_inv */ #(
            .INIT(32'b00000000000000100011111011001100))
        _N10183_1154_inv_vname (
            .Z (_N10183_1154_inv),
            .I0 (_N10183_3556),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1154_inv_vname.orig_name = _N10183_1154_inv;
	// LUT = (I1&~I3&~I4)|(~I1&I2&I3&~I4)|(ID&~I1&I3&~I4)|(I1&~I2&~I4)|(I0&~I1&~I2&~I3&I4) ;

    GTP_LUT5 /* _N10183_1169_inv */ #(
            .INIT(32'b00010111011101111111000111111111))
        _N10183_1169_inv_vname (
            .Z (_N10183_1169_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1169_inv_vname.orig_name = _N10183_1169_inv;
	// LUT = (~I3&~I4)|(I2&~I4)|(~I1&~I2&I4)|(~I0&~I2&I4)|(~I1&~I3)|(~I0&~I3)|(~I0&~I1) ;

    GTP_LUT5 /* _N10183_1172_inv */ #(
            .INIT(32'b00000101001001000010010011011111))
        _N10183_1172_inv_vname (
            .Z (_N10183_1172_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
    // defparam _N10183_1172_inv_vname.orig_name = _N10183_1172_inv;
	// LUT = (~I2&~I3&~I4)|(I1&~I3&~I4)|(~I0&~I3&~I4)|(I0&~I1&I2&I3&~I4)|(I0&~I1&I2&~I3&I4)|(~I0&~I2&I3&I4)|(~I0&I1&~I2) ;

    GTP_LUT5 /* _N10183_1188_inv */ #(
            .INIT(32'b00011100110100100100000011100110))
        _N10183_1188_inv_vname (
            .Z (_N10183_1188_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1188_inv_vname.orig_name = _N10183_1188_inv;
	// LUT = (I0&~I1&~I3&~I4)|(~I0&I1&~I3&~I4)|(~I0&I1&I2&~I4)|(I1&~I2&I3&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(I1&I2&~I3) ;

    GTP_LUT5 /* _N10183_1195_inv */ #(
            .INIT(32'b01111111011111110011011110110111))
        _N10183_1195_inv_vname (
            .Z (_N10183_1195_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1195_inv_vname.orig_name = _N10183_1195_inv;
	// LUT = (I0&I2&~I3&~I4)|(~I2&I4)|(~I0&I4)|(~I0&~I2)|(~I1) ;

    GTP_LUT5 /* _N10183_1204_inv */ #(
            .INIT(32'b01100110111111010011011011111101))
        _N10183_1204_inv_vname (
            .Z (_N10183_1204_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1204_inv_vname.orig_name = _N10183_1204_inv;
	// LUT = (~I1&I2&~I4)|(~I0&I1&I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(~I0&I1&~I2)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_1206_inv */ #(
            .INIT(32'b00000000110111110000000000000010))
        _N10183_1206_inv_vname (
            .Z (_N10183_1206_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1206_inv_vname.orig_name = _N10183_1206_inv;
	// LUT = (I1&~I3&I4)|(~I0&~I3&I4)|(I0&~I1&~I2&~I3) ;

    GTP_LUT5 /* _N10183_1241_inv */ #(
            .INIT(32'b01010111010001111100111111100111))
        _N10183_1241_inv_vname (
            .Z (_N10183_1241_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1241_inv_vname.orig_name = _N10183_1241_inv;
	// LUT = (I0&~I1&~I3&~I4)|(I1&I3&~I4)|(I1&I2&~I4)|(~I0&I3&I4)|(~I1&~I2)|(~I0&I1) ;

    GTP_LUT5M /* _N10183_1245_inv */ #(
            .INIT(32'b00000000000000100011111011001100))
        _N10183_1245_inv_vname (
            .Z (_N10183_1245_inv),
            .I0 (_N10183_3556),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1245_inv_vname.orig_name = _N10183_1245_inv;
	// LUT = (I1&~I3&~I4)|(~I1&I2&I3&~I4)|(ID&~I1&I3&~I4)|(I1&~I2&~I4)|(I0&~I1&~I2&~I3&I4) ;

    GTP_LUT5 /* _N10183_1260_inv */ #(
            .INIT(32'b00010111011101111111000111111111))
        _N10183_1260_inv_vname (
            .Z (_N10183_1260_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1260_inv_vname.orig_name = _N10183_1260_inv;
	// LUT = (~I3&~I4)|(I2&~I4)|(~I1&~I2&I4)|(~I0&~I2&I4)|(~I1&~I3)|(~I0&~I3)|(~I0&~I1) ;

    GTP_LUT5 /* _N10183_1263_inv */ #(
            .INIT(32'b00000101001001000010010011011111))
        _N10183_1263_inv_vname (
            .Z (_N10183_1263_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
    // defparam _N10183_1263_inv_vname.orig_name = _N10183_1263_inv;
	// LUT = (~I2&~I3&~I4)|(I1&~I3&~I4)|(~I0&~I3&~I4)|(I0&~I1&I2&I3&~I4)|(I0&~I1&I2&~I3&I4)|(~I0&~I2&I3&I4)|(~I0&I1&~I2) ;

    GTP_LUT5 /* _N10183_1279_inv */ #(
            .INIT(32'b00011100110100100100000011100110))
        _N10183_1279_inv_vname (
            .Z (_N10183_1279_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1279_inv_vname.orig_name = _N10183_1279_inv;
	// LUT = (I0&~I1&~I3&~I4)|(~I0&I1&~I3&~I4)|(~I0&I1&I2&~I4)|(I1&~I2&I3&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(I1&I2&~I3) ;

    GTP_LUT5 /* _N10183_1286_inv */ #(
            .INIT(32'b01111111011111110011011110110111))
        _N10183_1286_inv_vname (
            .Z (_N10183_1286_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1286_inv_vname.orig_name = _N10183_1286_inv;
	// LUT = (I0&I2&~I3&~I4)|(~I2&I4)|(~I0&I4)|(~I0&~I2)|(~I1) ;

    GTP_LUT5 /* _N10183_1295_inv */ #(
            .INIT(32'b01100110111111010011011011111101))
        _N10183_1295_inv_vname (
            .Z (_N10183_1295_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1295_inv_vname.orig_name = _N10183_1295_inv;
	// LUT = (~I1&I2&~I4)|(~I0&I1&I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(~I0&I1&~I2)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_1297_inv */ #(
            .INIT(32'b00000000110111110000000000000010))
        _N10183_1297_inv_vname (
            .Z (_N10183_1297_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1297_inv_vname.orig_name = _N10183_1297_inv;
	// LUT = (I1&~I3&I4)|(~I0&~I3&I4)|(I0&~I1&~I2&~I3) ;

    GTP_LUT5 /* _N10183_1332_inv */ #(
            .INIT(32'b01010111010001111100111111100111))
        _N10183_1332_inv_vname (
            .Z (_N10183_1332_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1332_inv_vname.orig_name = _N10183_1332_inv;
	// LUT = (I0&~I1&~I3&~I4)|(I1&I3&~I4)|(I1&I2&~I4)|(~I0&I3&I4)|(~I1&~I2)|(~I0&I1) ;

    GTP_LUT5M /* _N10183_1336_inv */ #(
            .INIT(32'b00000000000000100011111011001100))
        _N10183_1336_inv_vname (
            .Z (_N10183_1336_inv),
            .I0 (_N10183_3556),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1336_inv_vname.orig_name = _N10183_1336_inv;
	// LUT = (I1&~I3&~I4)|(~I1&I2&I3&~I4)|(ID&~I1&I3&~I4)|(I1&~I2&~I4)|(I0&~I1&~I2&~I3&I4) ;

    GTP_LUT5 /* _N10183_1351_inv */ #(
            .INIT(32'b00010111011101111111000111111111))
        _N10183_1351_inv_vname (
            .Z (_N10183_1351_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1351_inv_vname.orig_name = _N10183_1351_inv;
	// LUT = (~I3&~I4)|(I2&~I4)|(~I1&~I2&I4)|(~I0&~I2&I4)|(~I1&~I3)|(~I0&~I3)|(~I0&~I1) ;

    GTP_LUT5 /* _N10183_1354_inv */ #(
            .INIT(32'b00000101001001000010010011011111))
        _N10183_1354_inv_vname (
            .Z (_N10183_1354_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
    // defparam _N10183_1354_inv_vname.orig_name = _N10183_1354_inv;
	// LUT = (~I2&~I3&~I4)|(I1&~I3&~I4)|(~I0&~I3&~I4)|(I0&~I1&I2&I3&~I4)|(I0&~I1&I2&~I3&I4)|(~I0&~I2&I3&I4)|(~I0&I1&~I2) ;

    GTP_LUT5 /* _N10183_1370_inv */ #(
            .INIT(32'b00011100110100100100000011100110))
        _N10183_1370_inv_vname (
            .Z (_N10183_1370_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1370_inv_vname.orig_name = _N10183_1370_inv;
	// LUT = (I0&~I1&~I3&~I4)|(~I0&I1&~I3&~I4)|(~I0&I1&I2&~I4)|(I1&~I2&I3&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(I1&I2&~I3) ;

    GTP_LUT5 /* _N10183_1377_inv */ #(
            .INIT(32'b01111111011111110011011110110111))
        _N10183_1377_inv_vname (
            .Z (_N10183_1377_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1377_inv_vname.orig_name = _N10183_1377_inv;
	// LUT = (I0&I2&~I3&~I4)|(~I2&I4)|(~I0&I4)|(~I0&~I2)|(~I1) ;

    GTP_LUT5 /* _N10183_1386_inv */ #(
            .INIT(32'b01100110111111010011011011111101))
        _N10183_1386_inv_vname (
            .Z (_N10183_1386_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1386_inv_vname.orig_name = _N10183_1386_inv;
	// LUT = (~I1&I2&~I4)|(~I0&I1&I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(~I0&I1&~I2)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_1388_inv */ #(
            .INIT(32'b00000000110111110000000000000010))
        _N10183_1388_inv_vname (
            .Z (_N10183_1388_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1388_inv_vname.orig_name = _N10183_1388_inv;
	// LUT = (I1&~I3&I4)|(~I0&~I3&I4)|(I0&~I1&~I2&~I3) ;

    GTP_LUT5 /* _N10183_1423_inv */ #(
            .INIT(32'b01010111010001111100111111100111))
        _N10183_1423_inv_vname (
            .Z (_N10183_1423_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1423_inv_vname.orig_name = _N10183_1423_inv;
	// LUT = (I0&~I1&~I3&~I4)|(I1&I3&~I4)|(I1&I2&~I4)|(~I0&I3&I4)|(~I1&~I2)|(~I0&I1) ;

    GTP_LUT5M /* _N10183_1427_inv */ #(
            .INIT(32'b00000000000000100011111011001100))
        _N10183_1427_inv_vname (
            .Z (_N10183_1427_inv),
            .I0 (_N10183_3556),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1427_inv_vname.orig_name = _N10183_1427_inv;
	// LUT = (I1&~I3&~I4)|(~I1&I2&I3&~I4)|(ID&~I1&I3&~I4)|(I1&~I2&~I4)|(I0&~I1&~I2&~I3&I4) ;

    GTP_LUT5 /* _N10183_1442_inv */ #(
            .INIT(32'b00010111011101111111000111111111))
        _N10183_1442_inv_vname (
            .Z (_N10183_1442_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1442_inv_vname.orig_name = _N10183_1442_inv;
	// LUT = (~I3&~I4)|(I2&~I4)|(~I1&~I2&I4)|(~I0&~I2&I4)|(~I1&~I3)|(~I0&~I3)|(~I0&~I1) ;

    GTP_LUT5 /* _N10183_1445_inv */ #(
            .INIT(32'b00000101001001000010010011011111))
        _N10183_1445_inv_vname (
            .Z (_N10183_1445_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
    // defparam _N10183_1445_inv_vname.orig_name = _N10183_1445_inv;
	// LUT = (~I2&~I3&~I4)|(I1&~I3&~I4)|(~I0&~I3&~I4)|(I0&~I1&I2&I3&~I4)|(I0&~I1&I2&~I3&I4)|(~I0&~I2&I3&I4)|(~I0&I1&~I2) ;

    GTP_LUT5 /* _N10183_1461_inv */ #(
            .INIT(32'b00011100110100100100000011100110))
        _N10183_1461_inv_vname (
            .Z (_N10183_1461_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1461_inv_vname.orig_name = _N10183_1461_inv;
	// LUT = (I0&~I1&~I3&~I4)|(~I0&I1&~I3&~I4)|(~I0&I1&I2&~I4)|(I1&~I2&I3&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(I1&I2&~I3) ;

    GTP_LUT5 /* _N10183_1468_inv */ #(
            .INIT(32'b01111111011111110011011110110111))
        _N10183_1468_inv_vname (
            .Z (_N10183_1468_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1468_inv_vname.orig_name = _N10183_1468_inv;
	// LUT = (I0&I2&~I3&~I4)|(~I2&I4)|(~I0&I4)|(~I0&~I2)|(~I1) ;

    GTP_LUT5 /* _N10183_1477_inv */ #(
            .INIT(32'b01100110111111010011011011111101))
        _N10183_1477_inv_vname (
            .Z (_N10183_1477_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1477_inv_vname.orig_name = _N10183_1477_inv;
	// LUT = (~I1&I2&~I4)|(~I0&I1&I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(~I0&I1&~I2)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_1479_inv */ #(
            .INIT(32'b00000000110111110000000000000010))
        _N10183_1479_inv_vname (
            .Z (_N10183_1479_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1479_inv_vname.orig_name = _N10183_1479_inv;
	// LUT = (I1&~I3&I4)|(~I0&~I3&I4)|(I0&~I1&~I2&~I3) ;

    GTP_LUT5 /* _N10183_1514_inv */ #(
            .INIT(32'b01010111010001111100111111100111))
        _N10183_1514_inv_vname (
            .Z (_N10183_1514_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1514_inv_vname.orig_name = _N10183_1514_inv;
	// LUT = (I0&~I1&~I3&~I4)|(I1&I3&~I4)|(I1&I2&~I4)|(~I0&I3&I4)|(~I1&~I2)|(~I0&I1) ;

    GTP_LUT5M /* _N10183_1518_inv */ #(
            .INIT(32'b00000000000000100011111011001100))
        _N10183_1518_inv_vname (
            .Z (_N10183_1518_inv),
            .I0 (_N10183_3556),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1518_inv_vname.orig_name = _N10183_1518_inv;
	// LUT = (I1&~I3&~I4)|(~I1&I2&I3&~I4)|(ID&~I1&I3&~I4)|(I1&~I2&~I4)|(I0&~I1&~I2&~I3&I4) ;

    GTP_LUT5 /* _N10183_1533_inv */ #(
            .INIT(32'b00010111011101111111000111111111))
        _N10183_1533_inv_vname (
            .Z (_N10183_1533_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1533_inv_vname.orig_name = _N10183_1533_inv;
	// LUT = (~I3&~I4)|(I2&~I4)|(~I1&~I2&I4)|(~I0&~I2&I4)|(~I1&~I3)|(~I0&~I3)|(~I0&~I1) ;

    GTP_LUT5 /* _N10183_1536_inv */ #(
            .INIT(32'b00000101001001000010010011011111))
        _N10183_1536_inv_vname (
            .Z (_N10183_1536_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
    // defparam _N10183_1536_inv_vname.orig_name = _N10183_1536_inv;
	// LUT = (~I2&~I3&~I4)|(I1&~I3&~I4)|(~I0&~I3&~I4)|(I0&~I1&I2&I3&~I4)|(I0&~I1&I2&~I3&I4)|(~I0&~I2&I3&I4)|(~I0&I1&~I2) ;

    GTP_LUT5 /* _N10183_1552_inv */ #(
            .INIT(32'b00011100110100100100000011100110))
        _N10183_1552_inv_vname (
            .Z (_N10183_1552_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1552_inv_vname.orig_name = _N10183_1552_inv;
	// LUT = (I0&~I1&~I3&~I4)|(~I0&I1&~I3&~I4)|(~I0&I1&I2&~I4)|(I1&~I2&I3&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(I1&I2&~I3) ;

    GTP_LUT5 /* _N10183_1559_inv */ #(
            .INIT(32'b01111111011111110011011110110111))
        _N10183_1559_inv_vname (
            .Z (_N10183_1559_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1559_inv_vname.orig_name = _N10183_1559_inv;
	// LUT = (I0&I2&~I3&~I4)|(~I2&I4)|(~I0&I4)|(~I0&~I2)|(~I1) ;

    GTP_LUT5 /* _N10183_1568_inv */ #(
            .INIT(32'b01100110111111010011011011111101))
        _N10183_1568_inv_vname (
            .Z (_N10183_1568_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1568_inv_vname.orig_name = _N10183_1568_inv;
	// LUT = (~I1&I2&~I4)|(~I0&I1&I4)|(I1&~I3)|(~I0&~I3)|(I0&~I1&I3)|(~I0&I1&~I2)|(I0&~I1&I2) ;

    GTP_LUT5 /* _N10183_1570_inv */ #(
            .INIT(32'b00000000110111110000000000000010))
        _N10183_1570_inv_vname (
            .Z (_N10183_1570_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1570_inv_vname.orig_name = _N10183_1570_inv;
	// LUT = (I1&~I3&I4)|(~I0&~I3&I4)|(I0&~I1&~I2&~I3) ;

    GTP_LUT5 /* _N10183_1605_inv */ #(
            .INIT(32'b01010111010001111100111111100111))
        _N10183_1605_inv_vname (
            .Z (_N10183_1605_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1605_inv_vname.orig_name = _N10183_1605_inv;
	// LUT = (I0&~I1&~I3&~I4)|(I1&I3&~I4)|(I1&I2&~I4)|(~I0&I3&I4)|(~I1&~I2)|(~I0&I1) ;

    GTP_LUT5M /* _N10183_1609_inv */ #(
            .INIT(32'b00000000000000100011111011001100))
        _N10183_1609_inv_vname (
            .Z (_N10183_1609_inv),
            .I0 (_N10183_3556),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
    // defparam _N10183_1609_inv_vname.orig_name = _N10183_1609_inv;
	// LUT = (I1&~I3&~I4)|(~I1&I2&I3&~I4)|(ID&~I1&I3&~I4)|(I1&~I2&~I4)|(I0&~I1&~I2&~I3&I4) ;

    GTP_LUT5 /* _N10183_1624_inv */ #(
            .INIT(32'b00010111011101111111000111111111))
        _N10183_1624_inv_vname (
            .Z (_N10183_1624_inv),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
    // defparam _N10183_1624_inv_vname.orig_name = _N10183_1624_inv;
	// LUT = (~I3&~I4)|(I2&~I4)|(~I1&~I2&I4)|(~I0&~I2&I4)|(~I1&~I3)|(~I0&~I3)|(~I0&~I1) ;

(* PAP_IO_DIRECTION="OUTPUT", PAP_IO_LOC="J7", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUF /* lcd_bl_obuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        lcd_bl_obuf (
            .O (lcd_bl),
            .I (1'b1));
	// ../../rtl/top_lcd_touch.v:31

(* PAP_IO_DIRECTION="OUTPUT", PAP_IO_LOC="L5", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUF /* lcd_clk_obuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        lcd_clk_obuf (
            .O (lcd_clk),
            .I (nt_lcd_clk));
	// ../../rtl/top_lcd_touch.v:32

(* PAP_IO_DIRECTION="OUTPUT", PAP_IO_LOC="J6", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUF /* lcd_de_obuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        lcd_de_obuf (
            .O (lcd_de),
            .I (nt_lcd_de));
	// ../../rtl/top_lcd_touch.v:28

(* PAP_IO_DIRECTION="OUTPUT", PAP_IO_LOC="D1", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUF /* lcd_hs_obuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        lcd_hs_obuf (
            .O (lcd_hs),
            .I (1'b1));
	// ../../rtl/top_lcd_touch.v:29

(* PAP_IO_DIRECTION="OUTPUT", PAP_IO_LOC="F4", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUF /* lcd_rst_n_obuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        lcd_rst_n_obuf (
            .O (lcd_rst_n),
            .I (1'b1));
	// ../../rtl/top_lcd_touch.v:33

(* PAP_IO_DIRECTION="OUTPUT", PAP_IO_LOC="D2", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUF /* lcd_vs_obuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        lcd_vs_obuf (
            .O (lcd_vs),
            .I (1'b1));
	// ../../rtl/top_lcd_touch.v:30

(* PAP_IO_DIRECTION="INPUT", PAP_IO_LOC="V9", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_PULLUP="TRUE" *)    GTP_INBUF /* sys_clk_ibuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .TERM_DDR("ON"))
        sys_clk_ibuf (
            .O (nt_sys_clk),
            .I (sys_clk));
	// ../../rtl/top_lcd_touch.v:20

(* PAP_IO_DIRECTION="INPUT", PAP_IO_LOC="C4", PAP_IO_VCCIO="1.8", PAP_IO_STANDARD="LVCMOS18", PAP_IO_PULLUP="TRUE" *)    GTP_INBUF /* sys_rst_n_ibuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .TERM_DDR("ON"))
        sys_rst_n_ibuf (
            .O (nt_sys_rst_n),
            .I (sys_rst_n));
	// ../../rtl/top_lcd_touch.v:21

(* PAP_IO_DIRECTION="OUTPUT", PAP_IO_LOC="J1", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUF /* touch_rst_n_obuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        touch_rst_n_obuf (
            .O (touch_rst_n),
            .I (nt_touch_rst_n));
	// ../../rtl/top_lcd_touch.v:26

(* PAP_IO_DIRECTION="OUTPUT", PAP_IO_LOC="H6", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUF /* touch_scl_obuf */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        touch_scl_obuf (
            .O (touch_scl),
            .I (nt_touch_scl));
	// ../../rtl/top_lcd_touch.v:24

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="H3", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[0]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[0]  (
            .O (lcd_rgb[0]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="H4", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[1]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[1]  (
            .O (lcd_rgb[1]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="F1", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[2]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[2]  (
            .O (lcd_rgb[2]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="F2", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[3]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[3]  (
            .O (lcd_rgb[3]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="K1", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[4]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[4]  (
            .O (lcd_rgb[4]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="K2", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[5]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[5]  (
            .O (lcd_rgb[5]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="F5", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[6]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[6]  (
            .O (lcd_rgb[6]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="K5", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_IOBUF /* \u_lcd_rgb_char.lcd_rgb_tri[7]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"), 
            .TERM_DDR("ON"))
        \u_lcd_rgb_char.lcd_rgb_tri[7]  (
            .IO (lcd_rgb[7]),
            .O (_N0),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="E1", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[8]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[8]  (
            .O (lcd_rgb[8]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="E3", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[9]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[9]  (
            .O (lcd_rgb[9]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="L3", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[10]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[10]  (
            .O (lcd_rgb[10]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="L4", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[11]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[11]  (
            .O (lcd_rgb[11]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="K3", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[12]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[12]  (
            .O (lcd_rgb[12]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="K4", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[13]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[13]  (
            .O (lcd_rgb[13]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="K6", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[14]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[14]  (
            .O (lcd_rgb[14]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="L7", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_IOBUF /* \u_lcd_rgb_char.lcd_rgb_tri[15]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"), 
            .TERM_DDR("ON"))
        \u_lcd_rgb_char.lcd_rgb_tri[15]  (
            .IO (lcd_rgb[15]),
            .O (_N1),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="H1", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[16]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[16]  (
            .O (lcd_rgb[16]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="H2", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[17]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[17]  (
            .O (lcd_rgb[17]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="D3", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[18]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[18]  (
            .O (lcd_rgb[18]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="E4", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[19]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[19]  (
            .O (lcd_rgb[19]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="G6", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[20]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[20]  (
            .O (lcd_rgb[20]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="H7", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[21]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[21]  (
            .O (lcd_rgb[21]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="G1", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_lcd_rgb_char.lcd_rgb_tri[22]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_lcd_rgb_char.lcd_rgb_tri[22]  (
            .O (lcd_rgb[22]),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="G3", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_IOBUF /* \u_lcd_rgb_char.lcd_rgb_tri[23]  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"), 
            .TERM_DDR("ON"))
        \u_lcd_rgb_char.lcd_rgb_tri[23]  (
            .IO (lcd_rgb[23]),
            .O (_N2),
            .I (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .T (nt_lcd_de_inv));
	// ../../rtl/top_lcd_touch.v:34

    GTP_INV \u_lcd_rgb_char/u_binary2bcd_x/N0_vname  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .I (nt_sys_rst_n));
    // defparam \u_lcd_rgb_char/u_binary2bcd_x/N0_vname .orig_name = \u_lcd_rgb_char/u_binary2bcd_x/N0 ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N7_sum2  */ #(
            .INIT(8'b01101010))
        \u_lcd_rgb_char/u_binary2bcd_x/N7_sum2  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N7 [2] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [2] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [1] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [0] ));
	// LUT = (I0&~I2)|(~I0&I1&I2)|(I0&~I1) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_binary2bcd_x/N7_sum3  */ #(
            .INIT(16'b0110101010101010))
        \u_lcd_rgb_char/u_binary2bcd_x/N7_sum3  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N7 [3] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [3] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [2] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [1] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [0] ));
	// LUT = (I0&~I3)|(~I0&I1&I2&I3)|(I0&~I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N17_mux4_inv  */ #(
            .INIT(32'b01010101010101010101010101010111))
        \u_lcd_rgb_char/u_binary2bcd_x/N17_mux4_inv  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [4] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [3] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [1] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [0] ));
	// LUT = (~I1&~I2&~I3&~I4)|(~I0) ;

    GTP_LUT1 /* \u_lcd_rgb_char/u_binary2bcd_x/N19  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_binary2bcd_x/N19_vname  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N19 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
    // defparam \u_lcd_rgb_char/u_binary2bcd_x/N19_vname .orig_name = \u_lcd_rgb_char/u_binary2bcd_x/N19 ;
	// LUT = ~I0 ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_binary2bcd_x/N23_mux1  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_binary2bcd_x/N23_mux1  (
            .Z (_N48),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [17] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [16] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_binary2bcd_x/N23_mux3  */ #(
            .INIT(16'b1110111011101010))
        \u_lcd_rgb_char/u_binary2bcd_x/N23_mux3  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N23 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [19] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [18] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [17] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [16] ));
	// LUT = (I1&I3)|(I1&I2)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_binary2bcd_x/N31_mux1  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_binary2bcd_x/N31_mux1  (
            .Z (_N68),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [21] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [20] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_binary2bcd_x/N31_mux3  */ #(
            .INIT(16'b1110111011101010))
        \u_lcd_rgb_char/u_binary2bcd_x/N31_mux3  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N31 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [23] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [22] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [21] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [20] ));
	// LUT = (I1&I3)|(I1&I2)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_binary2bcd_x/N39_mux1  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_binary2bcd_x/N39_mux1  (
            .Z (_N88),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [25] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [24] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_binary2bcd_x/N39_mux3  */ #(
            .INIT(16'b1110111011101010))
        \u_lcd_rgb_char/u_binary2bcd_x/N39_mux3  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N39 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [27] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [26] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [25] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [24] ));
	// LUT = (I1&I3)|(I1&I2)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_binary2bcd_x/N47_mux1  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_binary2bcd_x/N47_mux1  (
            .Z (_N108),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [29] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [28] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_binary2bcd_x/N47_mux3  */ #(
            .INIT(16'b1110111011101010))
        \u_lcd_rgb_char/u_binary2bcd_x/N47_mux3  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N47 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [31] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [30] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [29] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [28] ));
	// LUT = (I1&I3)|(I1&I2)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N73_7  */ #(
            .INIT(32'b00000000000000100000000000000000))
        \u_lcd_rgb_char/u_binary2bcd_x/N73_7  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [4] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [3] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [1] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [0] ));
	// LUT = I0&~I1&~I2&~I3&I4 ;

    GTP_LUT1 /* \u_lcd_rgb_char/u_binary2bcd_x/N74  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_binary2bcd_x/N74  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N7 [0] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [0] ));
	// LUT = ~I0 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N76_1  */ #(
            .INIT(32'b00000000000000000000000000000001))
        \u_lcd_rgb_char/u_binary2bcd_x/N76_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [4] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [3] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [1] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [0] ));
	// LUT = ~I0&~I1&~I2&~I3&~I4 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N90[0]  */ #(
            .INIT(32'b00000000111111011111111100000000))
        \u_lcd_rgb_char/u_binary2bcd_x/N90[0]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N90 [1] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [4] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [3] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [1] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [0] ));
	// LUT = (I3&~I4)|(I2&~I3&I4)|(I1&~I3&I4)|(~I0&~I3&I4) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N90[1]  */ #(
            .INIT(32'b01101010101010001010101010101010))
        \u_lcd_rgb_char/u_binary2bcd_x/N90[1]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N90 [4] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [4] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [3] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [1] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [0] ));
	// LUT = (I0&~I4)|(~I0&I1&I2&I3&I4)|(I0&I1&~I3)|(I0&~I1&I3)|(I0&I1&~I2)|(I0&~I1&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_LUT2 /* \u_lcd_rgb_char/u_binary2bcd_x/N95  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_binary2bcd_x/N95_vname  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N95 ),
            .I0 (data[16]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
    // defparam \u_lcd_rgb_char/u_binary2bcd_x/N95_vname .orig_name = \u_lcd_rgb_char/u_binary2bcd_x/N95 ;
	// LUT = I0&I1 ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N97_1  */ #(
            .INIT(8'b11101010))
        \u_lcd_rgb_char/u_binary2bcd_x/N97_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
	// LUT = (I1&I2)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N98_7[0]_1  */ #(
            .INIT(32'b00000000110011000000000001011010))
        \u_lcd_rgb_char/u_binary2bcd_x/N98_7[0]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N98 [0] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [28] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [27] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N47 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
	// LUT = (I0&~I2&~I3&~I4)|(~I0&I2&~I3&~I4)|(I1&~I3&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N98_7[1]_1  */ #(
            .INIT(32'b00000000110011000000000010011010))
        \u_lcd_rgb_char/u_binary2bcd_x/N98_7[1]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N98 [1] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [29] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [28] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N47 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
	// LUT = (I0&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I1&~I3&I4)|(I0&I1&~I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_binary2bcd_x/N98_7[2]_1  */ #(
            .INIT(32'b00100010001000100000001000110000))
        \u_lcd_rgb_char/u_binary2bcd_x/N98_7[2]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N98 [2] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [29] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [30] ),
            .I3 (_N108),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .ID (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [31] ));
	// LUT = (~I1&I2&~I3&~I4)|(ID&~I1&~I2&I3&~I4)|(I0&~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N98_7[3]_1  */ #(
            .INIT(32'b00001100000001100000110000001010))
        \u_lcd_rgb_char/u_binary2bcd_x/N98_7[3]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N98 [3] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [31] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [30] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I4 (_N108));
	// LUT = (I0&I1&~I2&~I4)|(~I0&I1&~I2&I4)|(I0&~I1&~I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N104_7[0]_1  */ #(
            .INIT(32'b00000000110011000000000001011010))
        \u_lcd_rgb_char/u_binary2bcd_x/N104_7[0]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N104 [0] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [24] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [23] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N39 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
	// LUT = (I0&~I2&~I3&~I4)|(~I0&I2&~I3&~I4)|(I1&~I3&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N104_7[1]_1  */ #(
            .INIT(32'b00000000110011000000000010011010))
        \u_lcd_rgb_char/u_binary2bcd_x/N104_7[1]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N104 [1] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [25] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [24] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N39 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
	// LUT = (I0&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I1&~I3&I4)|(I0&I1&~I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_binary2bcd_x/N104_7[2]_1  */ #(
            .INIT(32'b00100010001000100000001000110000))
        \u_lcd_rgb_char/u_binary2bcd_x/N104_7[2]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N104 [2] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [25] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [26] ),
            .I3 (_N88),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .ID (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [27] ));
	// LUT = (~I1&I2&~I3&~I4)|(ID&~I1&~I2&I3&~I4)|(I0&~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N104_7[3]_1  */ #(
            .INIT(32'b00001100000001100000110000001010))
        \u_lcd_rgb_char/u_binary2bcd_x/N104_7[3]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N104 [3] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [27] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [26] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I4 (_N88));
	// LUT = (I0&I1&~I2&~I4)|(~I0&I1&~I2&I4)|(I0&~I1&~I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N110_7[0]_1  */ #(
            .INIT(32'b00000000110011000000000001011010))
        \u_lcd_rgb_char/u_binary2bcd_x/N110_7[0]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N110 [0] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [20] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [19] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N31 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
	// LUT = (I0&~I2&~I3&~I4)|(~I0&I2&~I3&~I4)|(I1&~I3&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N110_7[1]_1  */ #(
            .INIT(32'b00000000110011000000000010011010))
        \u_lcd_rgb_char/u_binary2bcd_x/N110_7[1]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N110 [1] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [21] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [20] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N31 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
	// LUT = (I0&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I1&~I3&I4)|(I0&I1&~I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_binary2bcd_x/N110_7[2]_1  */ #(
            .INIT(32'b00100010001000100000001000110000))
        \u_lcd_rgb_char/u_binary2bcd_x/N110_7[2]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N110 [2] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [21] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [22] ),
            .I3 (_N68),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .ID (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [23] ));
	// LUT = (~I1&I2&~I3&~I4)|(ID&~I1&~I2&I3&~I4)|(I0&~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N110_7[3]_1  */ #(
            .INIT(32'b00001100000001100000110000001010))
        \u_lcd_rgb_char/u_binary2bcd_x/N110_7[3]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N110 [3] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [23] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [22] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I4 (_N68));
	// LUT = (I0&I1&~I2&~I4)|(~I0&I1&~I2&I4)|(I0&~I1&~I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N116_7[0]_1  */ #(
            .INIT(32'b00000000110011000000000001011010))
        \u_lcd_rgb_char/u_binary2bcd_x/N116_7[0]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N116 [0] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [16] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [15] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N23 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
	// LUT = (I0&~I2&~I3&~I4)|(~I0&I2&~I3&~I4)|(I1&~I3&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N116_7[1]_1  */ #(
            .INIT(32'b00000000110011000000000010011010))
        \u_lcd_rgb_char/u_binary2bcd_x/N116_7[1]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N116 [1] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [17] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [16] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N23 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ));
	// LUT = (I0&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I1&~I3&I4)|(I0&I1&~I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_binary2bcd_x/N116_7[2]_1  */ #(
            .INIT(32'b00100010001000100000001000110000))
        \u_lcd_rgb_char/u_binary2bcd_x/N116_7[2]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N116 [2] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [17] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [18] ),
            .I3 (_N48),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .ID (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [19] ));
	// LUT = (~I1&I2&~I3&~I4)|(ID&~I1&~I2&I3&~I4)|(I0&~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_x/N116_7[3]_1  */ #(
            .INIT(32'b00001100000001100000110000001010))
        \u_lcd_rgb_char/u_binary2bcd_x/N116_7[3]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N116 [3] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [19] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [18] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I4 (_N48));
	// LUT = (I0&I1&~I2&~I4)|(~I0&I1&~I2&I4)|(I0&~I1&~I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[0]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[0]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [0] ),
            .I0 (data[17]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [0] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[1]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[1]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [1] ),
            .I0 (data[18]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [1] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[2]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[2]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [2] ),
            .I0 (data[19]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [2] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[3]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[3]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [3] ),
            .I0 (data[20]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [3] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[4]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[4]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [4] ),
            .I0 (data[21]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [4] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[5]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[5]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [5] ),
            .I0 (data[22]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [5] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[6]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[6]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [6] ),
            .I0 (data[23]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [6] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[7]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[7]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [7] ),
            .I0 (data[24]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [7] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[8]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[8]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [8] ),
            .I0 (data[25]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [8] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[9]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[9]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [9] ),
            .I0 (data[26]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [9] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[10]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[10]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [10] ),
            .I0 (data[27]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [10] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[11]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[11]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [11] ),
            .I0 (data[28]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [11] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[12]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[12]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [12] ),
            .I0 (data[29]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [12] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[13]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[13]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [13] ),
            .I0 (data[30]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [13] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_x/N122[14]  */ #(
            .INIT(8'b10101100))
        \u_lcd_rgb_char/u_binary2bcd_x/N122[14]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_x/N122 [14] ),
            .I0 (data[31]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [14] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_x/N76 ));
	// LUT = (I1&~I2)|(I0&I2) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[0]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [16] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[1]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [17] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[2]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [18] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[3]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [19] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[4]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [20] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[5]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [21] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[6]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [22] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[7]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [23] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[8]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [24] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[9]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [25] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[10]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [26] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[11]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [27] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[12]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [12] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [28] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[13]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [13] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [29] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[14]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [14] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [30] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/bcd_data[15]  (
            .Q (\u_lcd_rgb_char/bcd_data_x [15] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [31] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[0]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N7 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[1]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N90 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[2]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N7 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[3]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N7 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/cnt_shift[4]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/cnt_shift [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N90 [4] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[0]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N95 ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[1]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[2]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[3]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[4]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[5]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [4] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[6]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [5] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[7]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [6] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[8]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [7] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[9]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [8] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[10]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [9] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[11]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [10] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[12]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [12] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [11] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[13]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [13] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [12] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[14]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [14] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [13] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[15]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [15] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N122 [14] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[16]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[16]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [16] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N116 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[17]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[17]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [17] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N116 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[18]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[18]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [18] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N116 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[19]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[19]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [19] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N116 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[20]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[20]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [20] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N110 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[21]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[21]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [21] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N110 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[22]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[22]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [22] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N110 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[23]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[23]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [23] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N110 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[24]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[24]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [24] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N104 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[25]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[25]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [25] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N104 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[26]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[26]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [26] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N104 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[27]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[27]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [27] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N104 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[28]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[28]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [28] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N98 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[29]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[29]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [29] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N98 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[30]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[30]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [30] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N98 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_x/data_shift[31]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/data_shift[31]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/data_shift [31] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N98 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_C /* \u_lcd_rgb_char/u_binary2bcd_x/shift_flag  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_x/shift_flag_vname  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_x/N19 ));
    // defparam \u_lcd_rgb_char/u_binary2bcd_x/shift_flag_vname .orig_name = \u_lcd_rgb_char/u_binary2bcd_x/shift_flag ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:68

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N7_sum2  */ #(
            .INIT(8'b01111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N7_sum2  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N7 [2] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [0] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [1] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [2] ));
	// LUT = (I0&I1&~I2)|(~I1&I2)|(~I0&I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_binary2bcd_y/N7_sum3  */ #(
            .INIT(16'b0111111110000000))
        \u_lcd_rgb_char/u_binary2bcd_y/N7_sum3  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N7 [3] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [0] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [1] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [3] ));
	// LUT = (I0&I1&I2&~I3)|(~I2&I3)|(~I1&I3)|(~I0&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N17_mux4_inv  */ #(
            .INIT(32'b00000000000000011111111111111111))
        \u_lcd_rgb_char/u_binary2bcd_y/N17_mux4_inv  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [0] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [1] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [3] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [4] ));
	// LUT = (~I4)|(~I0&~I1&~I2&~I3) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_binary2bcd_y/N23_mux1  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_binary2bcd_y/N23_mux1  (
            .Z (_N154),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [16] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [17] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_binary2bcd_y/N23_mux3  */ #(
            .INIT(16'b1111111111100000))
        \u_lcd_rgb_char/u_binary2bcd_y/N23_mux3  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N23 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [16] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [17] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [18] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [19] ));
	// LUT = (I3)|(I1&I2)|(I0&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_binary2bcd_y/N31_mux1  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_binary2bcd_y/N31_mux1  (
            .Z (_N174),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [20] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [21] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_binary2bcd_y/N31_mux3  */ #(
            .INIT(16'b1111111111100000))
        \u_lcd_rgb_char/u_binary2bcd_y/N31_mux3  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N31 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [20] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [21] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [22] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [23] ));
	// LUT = (I3)|(I1&I2)|(I0&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_binary2bcd_y/N39_mux1  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_binary2bcd_y/N39_mux1  (
            .Z (_N194),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [24] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [25] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_binary2bcd_y/N39_mux3  */ #(
            .INIT(16'b1111111111100000))
        \u_lcd_rgb_char/u_binary2bcd_y/N39_mux3  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N39 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [24] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [25] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [26] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [27] ));
	// LUT = (I3)|(I1&I2)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N73_7  */ #(
            .INIT(32'b00000000000000100000000000000000))
        \u_lcd_rgb_char/u_binary2bcd_y/N73_7  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [0] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [1] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [3] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [4] ));
	// LUT = I0&~I1&~I2&~I3&I4 ;

    GTP_LUT1 /* \u_lcd_rgb_char/u_binary2bcd_y/N74  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_binary2bcd_y/N74  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N7 [0] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [0] ));
	// LUT = ~I0 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N76_1  */ #(
            .INIT(32'b00000000000000000000000000000001))
        \u_lcd_rgb_char/u_binary2bcd_y/N76_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [0] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [1] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [3] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [4] ));
	// LUT = ~I0&~I1&~I2&~I3&~I4 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N90[0]  */ #(
            .INIT(32'b01100110011001000110011001100110))
        \u_lcd_rgb_char/u_binary2bcd_y/N90[0]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N90 [1] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [0] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [1] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [3] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [4] ));
	// LUT = (I0&~I1&~I4)|(I0&~I1&I3)|(I0&~I1&I2)|(~I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N90[1]  */ #(
            .INIT(32'b01111111111111011000000000000000))
        \u_lcd_rgb_char/u_binary2bcd_y/N90[1]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N90 [4] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [0] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [1] ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [2] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [3] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [4] ));
	// LUT = (I0&I1&I2&I3&~I4)|(I1&~I3&I4)|(~I1&I3&I4)|(I1&~I2&I4)|(~I1&I2&I4)|(~I0&I4) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_LUT2 /* \u_lcd_rgb_char/u_binary2bcd_y/N95  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_binary2bcd_y/N95_vname  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N95 ),
            .I0 (data[0]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ));
    // defparam \u_lcd_rgb_char/u_binary2bcd_y/N95_vname .orig_name = \u_lcd_rgb_char/u_binary2bcd_y/N95 ;
	// LUT = I0&I1 ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N97_1  */ #(
            .INIT(8'b11101100))
        \u_lcd_rgb_char/u_binary2bcd_y/N97_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/N97 ));
	// LUT = (I0&I2)|(I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N104_7[0]_1  */ #(
            .INIT(32'b00001011000000010000111000000100))
        \u_lcd_rgb_char/u_binary2bcd_y/N104_7[0]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N104 [0] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N39 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [23] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [24] ));
	// LUT = (~I0&I1&~I2&~I4)|(~I0&~I1&~I2&I4)|(I0&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N104_7[1]_1  */ #(
            .INIT(32'b00001111000000010000101000000100))
        \u_lcd_rgb_char/u_binary2bcd_y/N104_7[1]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N104 [1] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N39 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [24] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [25] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&~I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_binary2bcd_y/N104_7[2]_1  */ #(
            .INIT(32'b00100010001000100001000000100010))
        \u_lcd_rgb_char/u_binary2bcd_y/N104_7[2]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N104 [2] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [25] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [27] ),
            .I3 (_N194),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .ID (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [26] ));
	// LUT = (ID&~I1&~I3&~I4)|(~ID&~I1&I2&I3&~I4)|(I0&~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N104_7[3]_1  */ #(
            .INIT(32'b00100001001100000011000100100000))
        \u_lcd_rgb_char/u_binary2bcd_y/N104_7[3]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N104 [3] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [26] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [27] ),
            .I4 (_N194));
	// LUT = (~I0&~I1&I3&~I4)|(~I1&I2&~I3&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N110_7[0]_1  */ #(
            .INIT(32'b00001011000000010000111000000100))
        \u_lcd_rgb_char/u_binary2bcd_y/N110_7[0]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N110 [0] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N31 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [19] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [20] ));
	// LUT = (~I0&I1&~I2&~I4)|(~I0&~I1&~I2&I4)|(I0&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N110_7[1]_1  */ #(
            .INIT(32'b00001111000000010000101000000100))
        \u_lcd_rgb_char/u_binary2bcd_y/N110_7[1]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N110 [1] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N31 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [20] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [21] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&~I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_binary2bcd_y/N110_7[2]_1  */ #(
            .INIT(32'b00100010001000100001000000100010))
        \u_lcd_rgb_char/u_binary2bcd_y/N110_7[2]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N110 [2] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [21] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [23] ),
            .I3 (_N174),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .ID (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [22] ));
	// LUT = (ID&~I1&~I3&~I4)|(~ID&~I1&I2&I3&~I4)|(I0&~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N110_7[3]_1  */ #(
            .INIT(32'b00100001001100000011000100100000))
        \u_lcd_rgb_char/u_binary2bcd_y/N110_7[3]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N110 [3] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [22] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [23] ),
            .I4 (_N174));
	// LUT = (~I0&~I1&I3&~I4)|(~I1&I2&~I3&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N116_7[0]_1  */ #(
            .INIT(32'b00001011000000010000111000000100))
        \u_lcd_rgb_char/u_binary2bcd_y/N116_7[0]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N116 [0] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N23 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [15] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [16] ));
	// LUT = (~I0&I1&~I2&~I4)|(~I0&~I1&~I2&I4)|(I0&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N116_7[1]_1  */ #(
            .INIT(32'b00001111000000010000101000000100))
        \u_lcd_rgb_char/u_binary2bcd_y/N116_7[1]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N116 [1] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N23 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [16] ),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [17] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&~I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_binary2bcd_y/N116_7[2]_1  */ #(
            .INIT(32'b00100010001000100001000000100010))
        \u_lcd_rgb_char/u_binary2bcd_y/N116_7[2]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N116 [2] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [17] ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [19] ),
            .I3 (_N154),
            .I4 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .ID (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [18] ));
	// LUT = (ID&~I1&~I3&~I4)|(~ID&~I1&I2&I3&~I4)|(I0&~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_binary2bcd_y/N116_7[3]_1  */ #(
            .INIT(32'b00100001001100000011000100100000))
        \u_lcd_rgb_char/u_binary2bcd_y/N116_7[3]_1  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N116 [3] ),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [18] ),
            .I3 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [19] ),
            .I4 (_N154));
	// LUT = (~I0&~I1&I3&~I4)|(~I1&I2&~I3&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[0]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[0]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [0] ),
            .I0 (data[1]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [0] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[1]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[1]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [1] ),
            .I0 (data[2]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [1] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[2]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[2]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [2] ),
            .I0 (data[3]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [2] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[3]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[3]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [3] ),
            .I0 (data[4]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [3] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[4]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[4]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [4] ),
            .I0 (data[5]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [4] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[5]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[5]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [5] ),
            .I0 (data[6]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [5] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[6]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[6]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [6] ),
            .I0 (data[7]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [6] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[7]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[7]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [7] ),
            .I0 (data[8]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [7] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[8]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[8]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [8] ),
            .I0 (data[9]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [8] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[9]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[9]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [9] ),
            .I0 (data[10]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [9] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[10]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[10]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [10] ),
            .I0 (data[11]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [10] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[11]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[11]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [11] ),
            .I0 (data[12]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [11] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[12]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[12]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [12] ),
            .I0 (data[13]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [12] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[13]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[13]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [13] ),
            .I0 (data[14]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [13] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT3 /* \u_lcd_rgb_char/u_binary2bcd_y/N122[14]  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_binary2bcd_y/N122[14]  (
            .Z (\u_lcd_rgb_char/u_binary2bcd_y/N122 [14] ),
            .I0 (data[15]),
            .I1 (\u_lcd_rgb_char/u_binary2bcd_y/N76 ),
            .I2 (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [14] ));
	// LUT = (~I1&I2)|(I0&I1) ;
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[0]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [16] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[1]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [17] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[2]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [18] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[3]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [19] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[4]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [20] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[5]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [21] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[6]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [22] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[7]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [23] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[8]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [24] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[9]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [25] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[10]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [26] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/bcd_data[11]  (
            .Q (\u_lcd_rgb_char/bcd_data_y [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N73 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [27] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:76

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[0]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N7 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[1]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N90 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[2]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N7 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[3]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N7 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/cnt_shift[4]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/cnt_shift [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N90 [4] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:38

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[0]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N95 ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[1]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[2]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[3]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[4]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[5]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [4] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[6]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [5] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[7]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [6] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[8]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [7] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[9]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [8] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[10]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [9] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[11]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [10] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[12]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [12] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [11] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[13]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [13] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [12] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[14]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [14] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [13] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[15]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [15] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N94 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N122 [14] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[16]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[16]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [16] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N116 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[17]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[17]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [17] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N116 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[18]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[18]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [18] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N116 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[19]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[19]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [19] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N116 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[20]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[20]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [20] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N110 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[21]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[21]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [21] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N110 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[22]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[22]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [22] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N110 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[23]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[23]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [23] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N110 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[24]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[24]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [24] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N104 [0] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[25]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[25]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [25] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N104 [1] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[26]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[26]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [26] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N104 [2] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_DFF_CE /* \u_lcd_rgb_char/u_binary2bcd_y/data_shift[27]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_binary2bcd_y/data_shift[27]  (
            .Q (\u_lcd_rgb_char/u_binary2bcd_y/data_shift [27] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_binary2bcd_y/N97 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_binary2bcd_y/N104 [3] ));
	// ../../rtl/lcd_rgb_char/binary2bcd.v:50

    GTP_LUT2 /* \u_lcd_rgb_char/u_clk_div/N19_1  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_clk_div/N19_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_clk_div/N19_2  */ #(
            .INIT(32'b01000010000000000000000000000000))
        \u_lcd_rgb_char/u_clk_div/N19_2  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I0 (lcd_id[8]),
            .I1 (lcd_id[12]),
            .I2 (lcd_id[13]),
            .I3 (_N10526),
            .I4 (_N10580));
	// LUT = (I0&~I1&~I2&I3&I4)|(~I0&I1&I2&I3&I4) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_clk_div/N33_7  */ #(
            .INIT(16'b0000001000000000))
        \u_lcd_rgb_char/u_clk_div/N33_7  (
            .Z (_N10584),
            .I0 (lcd_id[8]),
            .I1 (lcd_id[12]),
            .I2 (lcd_id[13]),
            .I3 (_N10526));
	// LUT = I0&~I1&~I2&I3 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_clk_div/N33_10  */ #(
            .INIT(32'b00000000001000000000000000000000))
        \u_lcd_rgb_char/u_clk_div/N33_10  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I0 (lcd_id[1]),
            .I1 (lcd_id[2]),
            .I2 (lcd_id[6]),
            .I3 (lcd_id[7]),
            .I4 (_N10584));
	// LUT = I0&~I1&I2&~I3&I4 ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_clk_div/N38_2  */ #(
            .INIT(8'b00100000))
        \u_lcd_rgb_char/u_clk_div/N38_2  (
            .Z (_N10585),
            .I0 (lcd_id[4]),
            .I1 (lcd_id[8]),
            .I2 (lcd_id[12]));
	// LUT = I0&~I1&I2 ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_clk_div/N39_1  */ #(
            .INIT(8'b00010000))
        \u_lcd_rgb_char/u_clk_div/N39_1  (
            .Z (_N10526),
            .I0 (lcd_id[3]),
            .I1 (lcd_id[4]),
            .I2 (lcd_id[14]));
	// LUT = ~I0&~I1&I2 ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_clk_div/N39_11  */ #(
            .INIT(16'b0000000000001000))
        \u_lcd_rgb_char/u_clk_div/N39_11  (
            .Z (_N11834),
            .I0 (lcd_id[1]),
            .I1 (lcd_id[2]),
            .I2 (lcd_id[6]),
            .I3 (lcd_id[7]));
	// LUT = I0&I1&~I2&~I3 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_clk_div/N39_13  */ #(
            .INIT(32'b01000000000000000000000000000000))
        \u_lcd_rgb_char/u_clk_div/N39_13  (
            .Z (\u_lcd_rgb_char/u_clk_div/N39 ),
            .I0 (lcd_id[3]),
            .I1 (lcd_id[13]),
            .I2 (lcd_id[14]),
            .I3 (_N10585),
            .I4 (_N11834));
	// LUT = ~I0&I1&I2&I3&I4 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_clk_div/N40  */ #(
            .INIT(32'b00000100000000000000000000000000))
        \u_lcd_rgb_char/u_clk_div/N40_vname  (
            .Z (\u_lcd_rgb_char/u_clk_div/N40 ),
            .I0 (lcd_id[1]),
            .I1 (lcd_id[2]),
            .I2 (lcd_id[6]),
            .I3 (lcd_id[7]),
            .I4 (_N10584));
    // defparam \u_lcd_rgb_char/u_clk_div/N40_vname .orig_name = \u_lcd_rgb_char/u_clk_div/N40 ;
	// LUT = ~I0&I1&~I2&I3&I4 ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_clk_div/N42_7  */ #(
            .INIT(16'b0000010000000000))
        \u_lcd_rgb_char/u_clk_div/N42_7  (
            .Z (_N10580),
            .I0 (lcd_id[1]),
            .I1 (lcd_id[2]),
            .I2 (lcd_id[6]),
            .I3 (lcd_id[7]));
	// LUT = ~I0&I1&~I2&I3 ;

    GTP_LUT1 /* \u_lcd_rgb_char/u_clk_div/N42_10_inv  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_clk_div/N42_10_inv  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb3 [8] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ));
	// LUT = ~I0 ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_clk_div/N42_14  */ #(
            .INIT(16'b0000000100000000))
        \u_lcd_rgb_char/u_clk_div/N42_14  (
            .Z (_N11824),
            .I0 (lcd_id[1]),
            .I1 (lcd_id[6]),
            .I2 (lcd_id[13]),
            .I3 (_N10585));
	// LUT = ~I0&~I1&~I2&I3 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_clk_div/N42_15  */ #(
            .INIT(32'b00000000000001000000000000000000))
        \u_lcd_rgb_char/u_clk_div/N42_15  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I0 (lcd_id[2]),
            .I1 (lcd_id[3]),
            .I2 (lcd_id[7]),
            .I3 (lcd_id[14]),
            .I4 (_N11824));
	// LUT = ~I0&I1&~I2&~I3&I4 ;

    GTP_DFF_CE /* \u_lcd_rgb_char/u_clk_div/clk_12_5m  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_clk_div/clk_12_5m_vname  (
            .Q (\u_lcd_rgb_char/u_clk_div/clk_12_5m ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (1'b1),
            .CLK (nt_sys_clk),
            .D (_N11805));
    // defparam \u_lcd_rgb_char/u_clk_div/clk_12_5m_vname .orig_name = \u_lcd_rgb_char/u_clk_div/clk_12_5m ;
	// ../../rtl/lcd_rgb_char/clk_div.v:43

    GTP_LUT2 /* \u_lcd_rgb_char/u_clk_div/clk_12_5m_ce_mux  */ #(
            .INIT(4'b0110))
        \u_lcd_rgb_char/u_clk_div/clk_12_5m_ce_mux  (
            .Z (_N11805),
            .I0 (\u_lcd_rgb_char/u_clk_div/clk_12_5m ),
            .I1 (\u_lcd_rgb_char/u_clk_div/div_4_cnt ));
	// LUT = I1^I0 ;

    GTP_DFF_C /* \u_lcd_rgb_char/u_clk_div/div_4_cnt  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_clk_div/div_4_cnt_vname  (
            .Q (\u_lcd_rgb_char/u_clk_div/div_4_cnt ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_clk_div/N3 ));
    // defparam \u_lcd_rgb_char/u_clk_div/div_4_cnt_vname .orig_name = \u_lcd_rgb_char/u_clk_div/div_4_cnt ;
	// ../../rtl/lcd_rgb_char/clk_div.v:43

    GTP_LUT1 /* \u_lcd_rgb_char/u_clk_div/div_4_cnt_inv  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_clk_div/div_4_cnt_inv  (
            .Z (\u_lcd_rgb_char/u_clk_div/N3 ),
            .I0 (\u_lcd_rgb_char/u_clk_div/div_4_cnt ));
	// LUT = ~I0 ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_clk_div/lcd_pclk_or[0]_2  */ #(
            .INIT(16'b1110101011000000))
        \u_lcd_rgb_char/u_clk_div/lcd_pclk_or[0]_2  (
            .Z (_N11839),
            .I0 (\u_lcd_rgb_char/u_binary2bcd_x/shift_flag ),
            .I1 (\u_lcd_rgb_char/u_clk_div/clk_12_5m ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ));
	// LUT = (I0&I3)|(I1&I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_clk_div/lcd_pclk_or[0]_3  */ #(
            .INIT(16'b1111111110101000))
        \u_lcd_rgb_char/u_clk_div/lcd_pclk_or[0]_3  (
            .Z (nt_lcd_clk),
            .I0 (nt_sys_clk),
            .I1 (\u_lcd_rgb_char/u_clk_div/N39 ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I3 (_N11839));
	// LUT = (I3)|(I0&I2)|(I0&I1) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_0  */ #(
            .INIT(32'b00110011001100110000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [0] ),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [1] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = ~I1 ;
	// CARRY = (1'b0) ? CIN : (~I1) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_1  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [1] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [6] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [0] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [2] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_2  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [2] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [7] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [1] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [3] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_3  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [3] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [8] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [2] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [4] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_4  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [4] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [9] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [3] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [5] ),
            .I2 (),
            .I3 (),
            .I4 (1'b1),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_5  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_5  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [5] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [10] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [4] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [6] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_6  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_6  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [6] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [11] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [5] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [7] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_7  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_7  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [7] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [12] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [6] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [8] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_8  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_8  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [8] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [13] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [7] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [9] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_9  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_9  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N46_1.co [9] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [14] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [8] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [10] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_10  */ #(
            .INIT(32'b01010101010101011111111111111111), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N46_1.fsub_10  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_display/N392 [15] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N46_1.co [9] ),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~CIN ;
	// CARRY = (1'b1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_0  */ #(
            .INIT(32'b00000000000000000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [0] ),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = (1'b0) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_1  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [1] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [0] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w[0]_inv ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/pixel_ypos_w[0]_inv ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_2  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [2] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [1] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [1] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/pixel_ypos_w [1] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_3  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [3] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [2] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [6] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [6] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_4  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [4] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [3] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [7] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [7] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_5  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_5  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [5] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [4] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [8] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [8] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_6  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_6  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [6] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [9] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [5] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [9] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [9] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_7  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_7  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [7] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [10] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [6] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [10] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [10] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_8  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_8  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [8] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [11] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [7] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [11] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [11] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_9  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_9  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [9] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [12] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [8] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [12] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [12] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_10  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_10  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [10] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [13] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [9] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [13] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [13] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_11  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_11  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [11] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [14] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [10] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [14] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [14] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_12  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_12  (
            .COUT (\u_lcd_rgb_char/u_lcd_display/N59_1.co [12] ),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [15] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [11] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [15] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [15] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_13  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_display/N59_1.fsub_13  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_display/N59 [16] ),
            .CIN (\u_lcd_rgb_char/u_lcd_display/N59_1.co [12] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N392 [15] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N392 [15] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_display.v:123

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_4570_4  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4570_4  (
            .Z (_N12187),
            .I0 (\u_lcd_rgb_char/pixel_ypos_w [6] ),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [7] ),
            .I2 (\u_lcd_rgb_char/pixel_ypos_w [10] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4570_6  */ #(
            .INIT(32'b11111111111111111111111011111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4570_6  (
            .Z (_N12189),
            .I0 (\u_lcd_rgb_char/pixel_ypos_w [5] ),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [8] ),
            .I2 (\u_lcd_rgb_char/pixel_ypos_w [9] ),
            .I3 (_N10183_31),
            .I4 (_N12187));
	// LUT = (I4)|(~I0&~I3)|(I0&I3)|(I2)|(I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4570_8  */ #(
            .INIT(32'b11111111111010101111111111101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4570_8  (
            .Z (\u_lcd_rgb_char/u_lcd_display/N9971 [0] ),
            .I0 (_N10183_6),
            .I1 (_N10183_5),
            .I2 (_N10183_9),
            .I3 (_N12189),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [5] ),
            .ID (_N10183_7));
	// LUT = (ID&~I4)|(I0&I4)|(I3)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4574_4  */ #(
            .INIT(32'b11111111111111111111111110011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4574_4  (
            .Z (_N10183_5),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .I2 (_N10183_20),
            .I3 (_N10183_36),
            .I4 (_N10183_62));
	// LUT = (I4)|(I3)|(~I2)|(~I0&~I1)|(I0&I1) ;

    GTP_MUX2LUT8 \u_lcd_rgb_char/u_lcd_display/N9971_4575  (
            .Z (_N10183_6),
            .I0 (_N10183_12),
            .I1 (_N10183_11),
            .S (\u_lcd_rgb_char/pixel_xpos_w [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4576  */ #(
            .INIT(32'b10101010111100000000000000100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4576  (
            .Z (_N10183_7),
            .I0 (_N10183_25),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .I2 (_N10183_26),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [4] ),
            .ID (_N10183_28));
	// LUT = (ID&~I1&~I3&~I4)|(I2&~I3&I4)|(I0&I3&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4578  (
            .Z (_N10183_9),
            .I0 (_N10183_17),
            .I1 (_N10183_18),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4580  (
            .Z (_N10183_11),
            .I0 (_N10183_22),
            .I1 (_N10183_21),
            .S (\u_lcd_rgb_char/pixel_xpos_w [6] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4581  (
            .Z (_N10183_12),
            .I0 (_N10183_24),
            .I1 (_N10183_23),
            .S (\u_lcd_rgb_char/pixel_xpos_w [6] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4586  */ #(
            .INIT(32'b11111111101010101111111111100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4586  (
            .Z (_N10183_17),
            .I0 (_N10183_58),
            .I1 (_N10183_62),
            .I2 (_N10183_97),
            .I3 (_N10183_36),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_98));
	// LUT = (I1&I2&~I4)|(ID&~I1&~I4)|(I0&I4)|(I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4587  */ #(
            .INIT(32'b11111111111111101110111011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4587  (
            .Z (_N10183_18),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (_N10183_36),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I3 (_N10183_172),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (_N10183_59));
	// LUT = (ID&~I4)|(I3&I4)|(I2&I4)|(I0&I4)|(I1) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_4589_6  */ #(
            .INIT(16'b1111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4589_6  (
            .Z (_N11868),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [9] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [10] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [12] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4589_8  */ #(
            .INIT(32'b11111111111111111111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4589_8  (
            .Z (_N10183_20),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [13] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [14] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [16] ),
            .I4 (_N11868));
	// LUT = (I4)|(I3)|(I2)|(I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4590  (
            .Z (_N10183_21),
            .I0 (_N10183_41),
            .I1 (_N10183_40),
            .S (\u_lcd_rgb_char/pixel_xpos_w [3] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4591  (
            .Z (_N10183_22),
            .I0 (_N10183_43),
            .I1 (_N10183_42),
            .S (\u_lcd_rgb_char/pixel_xpos_w [3] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4592  (
            .Z (_N10183_23),
            .I0 (_N10183_45),
            .I1 (_N10183_44),
            .S (\u_lcd_rgb_char/pixel_xpos_w [3] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4593  (
            .Z (_N10183_24),
            .I0 (_N10183_47),
            .I1 (_N10183_46),
            .S (\u_lcd_rgb_char/pixel_xpos_w [3] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4594  (
            .Z (_N10183_25),
            .I0 (_N10183_49),
            .I1 (_N10183_48),
            .S (\u_lcd_rgb_char/pixel_xpos_w [3] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4595  (
            .Z (_N10183_26),
            .I0 (_N10183_51),
            .I1 (_N10183_50),
            .S (\u_lcd_rgb_char/pixel_xpos_w [3] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4597  (
            .Z (_N10183_28),
            .I0 (_N10183_53),
            .I1 (_N10183_52),
            .S (\u_lcd_rgb_char/pixel_xpos_w [3] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4600_5  */ #(
            .INIT(32'b11111111111111111111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4600_5  (
            .Z (_N10183_31),
            .I0 (\u_lcd_rgb_char/pixel_ypos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_ypos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_ypos_w [2] ),
            .I3 (\u_lcd_rgb_char/pixel_ypos_w [3] ),
            .I4 (\u_lcd_rgb_char/pixel_ypos_w [4] ));
	// LUT = (I4)|(I3)|(I2)|(I1)|(I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_4605_3  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4605_3  (
            .Z (_N10183_36),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [8] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [10] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4609  */ #(
            .INIT(32'b11111010110110000111001001010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4609  (
            .Z (_N10183_40),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_69),
            .I3 (_N10183_104),
            .I4 (_N10183_105));
	// LUT = (I0&I1&I4)|(I0&~I1&I3)|(~I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4610  */ #(
            .INIT(32'b11001111010001111000101100000011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4610  (
            .Z (_N10183_41),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I2 (_N10183_71),
            .I3 (_N10183_108),
            .I4 (_N10183_109));
	// LUT = (~I0&I1&I4)|(I0&I1&I3)|(~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4611  */ #(
            .INIT(32'b11111010110110000111001001010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4611  (
            .Z (_N10183_42),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_73),
            .I3 (_N10183_112),
            .I4 (_N10183_113));
	// LUT = (I0&I1&I4)|(I0&~I1&I3)|(~I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4612  */ #(
            .INIT(32'b11001111010001111000101100000011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4612  (
            .Z (_N10183_43),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I2 (_N10183_75),
            .I3 (_N10183_116),
            .I4 (_N10183_117));
	// LUT = (~I0&I1&I4)|(I0&I1&I3)|(~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4613  */ #(
            .INIT(32'b11111010110110000111001001010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4613  (
            .Z (_N10183_44),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_77),
            .I3 (_N10183_120),
            .I4 (_N10183_121));
	// LUT = (I0&I1&I4)|(I0&~I1&I3)|(~I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4614  */ #(
            .INIT(32'b11001111010001111000101100000011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4614  (
            .Z (_N10183_45),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I2 (_N10183_79),
            .I3 (_N10183_124),
            .I4 (_N10183_125));
	// LUT = (~I0&I1&I4)|(I0&I1&I3)|(~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4615  */ #(
            .INIT(32'b11111010110110000111001001010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4615  (
            .Z (_N10183_46),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_81),
            .I3 (_N10183_128),
            .I4 (_N10183_129));
	// LUT = (I0&I1&I4)|(I0&~I1&I3)|(~I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4616  */ #(
            .INIT(32'b11001111010001111000101100000011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4616  (
            .Z (_N10183_47),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I2 (_N10183_83),
            .I3 (_N10183_132),
            .I4 (_N10183_133));
	// LUT = (~I0&I1&I4)|(I0&I1&I3)|(~I1&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4617  (
            .Z (_N10183_48),
            .I0 (_N10183_85),
            .I1 (_N10183_84),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4618  (
            .Z (_N10183_49),
            .I0 (_N10183_87_inv),
            .I1 (_N10183_86),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4619  (
            .Z (_N10183_50),
            .I0 (_N10183_89),
            .I1 (_N10183_88),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4620  (
            .Z (_N10183_51),
            .I0 (_N10183_91_inv),
            .I1 (_N10183_90),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4621  (
            .Z (_N10183_52),
            .I0 (_N10183_93),
            .I1 (_N10183_92),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4622  (
            .Z (_N10183_53),
            .I0 (_N10183_95_inv),
            .I1 (_N10183_94),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4627  */ #(
            .INIT(32'b11111111101010101110001011100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4627  (
            .Z (_N10183_58),
            .I0 (_N11364_2),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_167),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .I4 (_N10183_62),
            .ID (_N10183_166));
	// LUT = (I1&I2&~I4)|(ID&~I1&~I4)|(I3&I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4628  (
            .Z (_N10183_59),
            .I0 (_N10183_102),
            .I1 (_N10183_101),
            .S (_N10183_62));

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_4631  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4631  (
            .Z (_N10183_62),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [4] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [5] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4638  */ #(
            .INIT(32'b11011101110110000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4638  (
            .Z (_N10183_69),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (_N10183_180),
            .I2 (_N10183_317),
            .I3 (_N10183_318),
            .I4 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .ID (_N10183_106));
	// LUT = (~ID&~I4)|(~I0&I3&I4)|(~I0&I2&I4)|(I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4640  */ #(
            .INIT(32'b11101110001000100001110100011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4640  (
            .Z (_N10183_71),
            .I0 (_N10183_186),
            .I1 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I2 (_N10183_187),
            .I3 (_N10183_188),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (_N10183_185));
	// LUT = (I1&~I2&~I4)|(~ID&~I1&~I4)|(I1&I3&I4)|(I0&~I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4642  */ #(
            .INIT(32'b11011101110110000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4642  (
            .Z (_N10183_73),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (_N10183_196),
            .I2 (_N10183_317),
            .I3 (_N10183_349),
            .I4 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .ID (_N10183_114));
	// LUT = (~ID&~I4)|(~I0&I3&I4)|(~I0&I2&I4)|(I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4644  */ #(
            .INIT(32'b11101110001000100001110100011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4644  (
            .Z (_N10183_75),
            .I0 (_N10183_202),
            .I1 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I2 (_N10183_203),
            .I3 (_N10183_204),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (_N10183_201));
	// LUT = (I1&~I2&~I4)|(~ID&~I1&~I4)|(I1&I3&I4)|(I0&~I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4646  */ #(
            .INIT(32'b11011101110110000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4646  (
            .Z (_N10183_77),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (_N10183_212),
            .I2 (_N10183_317),
            .I3 (_N10183_380),
            .I4 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .ID (_N10183_122));
	// LUT = (~ID&~I4)|(~I0&I3&I4)|(~I0&I2&I4)|(I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4648  */ #(
            .INIT(32'b11101110001000100001110100011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4648  (
            .Z (_N10183_79),
            .I0 (_N10183_218),
            .I1 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I2 (_N10183_219),
            .I3 (_N10183_220),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (_N10183_217));
	// LUT = (I1&~I2&~I4)|(~ID&~I1&~I4)|(I1&I3&I4)|(I0&~I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4650  */ #(
            .INIT(32'b11011101110110000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4650  (
            .Z (_N10183_81),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (_N10183_228),
            .I2 (_N10183_317),
            .I3 (_N10183_411),
            .I4 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .ID (_N10183_130));
	// LUT = (~ID&~I4)|(~I0&I3&I4)|(~I0&I2&I4)|(I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4652  */ #(
            .INIT(32'b11101110001000100001110100011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4652  (
            .Z (_N10183_83),
            .I0 (_N10183_234),
            .I1 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I2 (_N10183_235),
            .I3 (_N10183_236),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (_N10183_233));
	// LUT = (I1&~I2&~I4)|(~ID&~I1&~I4)|(I1&I3&I4)|(I0&~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4653  */ #(
            .INIT(32'b11110011110100011110001011000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4653  (
            .Z (_N10183_84),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_137),
            .I3 (_N10183_237),
            .I4 (_N10183_238));
	// LUT = (~I0&~I1&I4)|(I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4654  */ #(
            .INIT(32'b11011101110110000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4654  (
            .Z (_N10183_85),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (_N10183_244),
            .I2 (_N10183_317),
            .I3 (_N10183_442),
            .I4 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .ID (_N10183_138));
	// LUT = (~ID&~I4)|(~I0&I3&I4)|(~I0&I2&I4)|(I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4655  */ #(
            .INIT(32'b10101010101010101101110111011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4655  (
            .Z (_N10183_86),
            .I0 (_N10183_140),
            .I1 (_N10183_248),
            .I2 (_N10183_449),
            .I3 (_N10183_450),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~ID&I3&~I4)|(~ID&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4657  */ #(
            .INIT(32'b11110011110100011110001011000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4657  (
            .Z (_N10183_88),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_145),
            .I3 (_N10183_253),
            .I4 (_N10183_254));
	// LUT = (~I0&~I1&I4)|(I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4658  */ #(
            .INIT(32'b11011101110110000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4658  (
            .Z (_N10183_89),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (_N10183_260),
            .I2 (_N10183_317),
            .I3 (_N10183_473),
            .I4 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .ID (_N10183_146));
	// LUT = (~ID&~I4)|(~I0&I3&I4)|(~I0&I2&I4)|(I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4659  */ #(
            .INIT(32'b10101010101010101101110111011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4659  (
            .Z (_N10183_90),
            .I0 (_N10183_148),
            .I1 (_N10183_264),
            .I2 (_N10183_480),
            .I3 (_N10183_481),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~ID&I3&~I4)|(~ID&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4661  */ #(
            .INIT(32'b11110011110100011110001011000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4661  (
            .Z (_N10183_92),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_153),
            .I3 (_N10183_269),
            .I4 (_N10183_270));
	// LUT = (~I0&~I1&I4)|(I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4662  */ #(
            .INIT(32'b11011101110110000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4662  (
            .Z (_N10183_93),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (_N10183_276),
            .I2 (_N10183_317),
            .I3 (_N10183_504),
            .I4 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .ID (_N10183_154));
	// LUT = (~ID&~I4)|(~I0&I3&I4)|(~I0&I2&I4)|(I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4663  */ #(
            .INIT(32'b10101010101010101101110111011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4663  (
            .Z (_N10183_94),
            .I0 (_N10183_156),
            .I1 (_N10183_280),
            .I2 (_N10183_511),
            .I3 (_N10183_512),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~ID&I3&~I4)|(~ID&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_4666  */ #(
            .INIT(16'b1111000111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4666  (
            .Z (_N10183_97),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_160),
            .I3 (_N10183_286));
	// LUT = (I0&~I3)|(I2)|(~I0&~I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4667  (
            .Z (_N10183_98),
            .I0 (_N10183_162),
            .I1 (_N10183_163),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4670  */ #(
            .INIT(32'b11111100101011001111110010101100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4670  (
            .Z (_N10183_101),
            .I0 (_N10183_543),
            .I1 (_N10183_168),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (_N10183_542));
	// LUT = (ID&I2&~I4)|(I0&I2&I4)|(I2&I3)|(I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4671  */ #(
            .INIT(32'b10101010101010101110111011100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4671  (
            .Z (_N10183_102),
            .I0 (_N10183_171),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I3 (_N10183_544),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .ID (_N10183_300));
	// LUT = (I1&I3&~I4)|(I1&I2&~I4)|(ID&~I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4673  */ #(
            .INIT(32'b11011111000100001110111100100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4673  (
            .Z (_N10183_104),
            .I0 (_N10183_554),
            .I1 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N12317),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_555));
	// LUT = (ID&~I1&I2&~I4)|(~I0&~I1&I2&I4)|(~I2&I3)|(I1&I3) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4674  (
            .Z (_N10183_105),
            .I0 (_N10183_175),
            .I1 (_N10183_176),
            .S (\u_lcd_rgb_char/bcd_data_y [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4675  (
            .Z (_N10183_106),
            .I0 (_N10183_178),
            .I1 (_N10183_177),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4677  (
            .Z (_N10183_108),
            .I0 (_N10183_181),
            .I1 (_N10183_182),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4678  */ #(
            .INIT(32'b11111111000011111111101100001011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4678  (
            .Z (_N10183_109),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_184),
            .I4 (_N10183_325));
	// LUT = (~I2&I4)|(I2&I3)|(~I1&~I2)|(I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4681  (
            .Z (_N10183_112),
            .I0 (_N10183_190),
            .I1 (_N10183_189),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4682  (
            .Z (_N10183_113),
            .I0 (_N10183_191),
            .I1 (_N10183_192),
            .S (\u_lcd_rgb_char/bcd_data_x [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4683  (
            .Z (_N10183_114),
            .I0 (_N10183_194),
            .I1 (_N10183_193),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4685  (
            .Z (_N10183_116),
            .I0 (_N10183_197),
            .I1 (_N10183_198),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4686  */ #(
            .INIT(32'b11111111000011111111101100001011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4686  (
            .Z (_N10183_117),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_200),
            .I4 (_N10183_356));
	// LUT = (~I2&I4)|(I2&I3)|(~I1&~I2)|(I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4689  (
            .Z (_N10183_120),
            .I0 (_N10183_206),
            .I1 (_N10183_205),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4690  (
            .Z (_N10183_121),
            .I0 (_N10183_207),
            .I1 (_N10183_208),
            .S (\u_lcd_rgb_char/bcd_data_y [6] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4691  (
            .Z (_N10183_122),
            .I0 (_N10183_210),
            .I1 (_N10183_209),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4693  (
            .Z (_N10183_124),
            .I0 (_N10183_213),
            .I1 (_N10183_214),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4694  */ #(
            .INIT(32'b11111111000011111111101100001011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4694  (
            .Z (_N10183_125),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_216),
            .I4 (_N10183_387));
	// LUT = (~I2&I4)|(I2&I3)|(~I1&~I2)|(I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4697  (
            .Z (_N10183_128),
            .I0 (_N10183_222),
            .I1 (_N10183_221),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4698  (
            .Z (_N10183_129),
            .I0 (_N10183_223),
            .I1 (_N10183_224),
            .S (\u_lcd_rgb_char/bcd_data_x [6] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4699  (
            .Z (_N10183_130),
            .I0 (_N10183_226),
            .I1 (_N10183_225),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4701  (
            .Z (_N10183_132),
            .I0 (_N10183_229),
            .I1 (_N10183_230),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4702  */ #(
            .INIT(32'b11111111000011111111101100001011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4702  (
            .Z (_N10183_133),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_232),
            .I4 (_N10183_418));
	// LUT = (~I2&I4)|(I2&I3)|(~I1&~I2)|(I0&~I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4706  (
            .Z (_N10183_137),
            .I0 (_N10183_239),
            .I1 (_N10183_240),
            .S (\u_lcd_rgb_char/bcd_data_y [10] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4707  (
            .Z (_N10183_138),
            .I0 (_N10183_242),
            .I1 (_N10183_241),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4709  (
            .Z (_N10183_140),
            .I0 (_N10183_245),
            .I1 (_N10183_246),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4714  (
            .Z (_N10183_145),
            .I0 (_N10183_255),
            .I1 (_N10183_256),
            .S (\u_lcd_rgb_char/bcd_data_x [10] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4715  (
            .Z (_N10183_146),
            .I0 (_N10183_258),
            .I1 (_N10183_257),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4717  (
            .Z (_N10183_148),
            .I0 (_N10183_261),
            .I1 (_N10183_262),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4722  (
            .Z (_N10183_153),
            .I0 (_N10183_271),
            .I1 (_N10183_272),
            .S (\u_lcd_rgb_char/bcd_data_x [14] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4723  (
            .Z (_N10183_154),
            .I0 (_N10183_274),
            .I1 (_N10183_273),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4725  (
            .Z (_N10183_156),
            .I0 (_N10183_277),
            .I1 (_N10183_278),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_4729  */ #(
            .INIT(16'b1111111100000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_4729  (
            .Z (_N10183_160),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [7] ));
	// LUT = (I3)|(~I0&~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4731  */ #(
            .INIT(32'b11111111111100001101111111010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4731  (
            .Z (_N10183_162),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .I3 (_N10183_288),
            .I4 (_N10183_527));
	// LUT = (I2&I4)|(~I2&I3)|(I1&I2)|(~I0&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4732  */ #(
            .INIT(32'b11111111011111101010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4732  (
            .Z (_N10183_163),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (_N11860),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .ID (_N10183_290));
	// LUT = (ID&~I4)|(I3&I4)|(I0&~I2&I4)|(~I0&I2&I4)|(I0&~I1&I4)|(~I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4735  */ #(
            .INIT(32'b11100010111111111110001011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4735  (
            .Z (_N10183_166),
            .I0 (_N10183_964),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .I2 (_N10183_535),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .ID (_N10183_292));
	// LUT = (ID&~I1&~I4)|(I0&~I1&I4)|(~I3)|(I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4736  (
            .Z (_N10183_167),
            .I0 (_N10183_296),
            .I1 (_N10183_295),
            .S (\u_lcd_rgb_char/pixel_xpos_w [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4737  */ #(
            .INIT(32'b11111111111111110001000000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4737  (
            .Z (_N10183_168),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I4 (_N10183_160));
	// LUT = (I4)|(~I0&~I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4740  (
            .Z (_N10183_171),
            .I0 (_N10183_301),
            .I1 (_N10183_302),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4741  */ #(
            .INIT(32'b11111111110010101111101011001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4741  (
            .Z (_N10183_172),
            .I0 (_N10183_983),
            .I1 (_N10183_551),
            .I2 (_N10183_62),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .ID (_N10924_2));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(I0&~I2&I4)|(I2&I3)|(ID&I3)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4743  */ #(
            .INIT(32'b11111100101110000111010000110000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4743  (
            .Z (_N10183_174),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_307),
            .I3 (_N10183_560),
            .I4 (_N10183_561));
	// LUT = (I0&I1&I4)|(~I0&I1&I3)|(~I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4744  (
            .Z (_N10183_175),
            .I0 (_N10183_310),
            .I1 (_N10183_309),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4745  (
            .Z (_N10183_176),
            .I0 (_N10183_311),
            .I1 (_N10183_312),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4746  */ #(
            .INIT(32'b10100000101000110101001101010011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4746  (
            .Z (_N10183_177),
            .I0 (_N10183_572),
            .I1 (_N10183_571),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_573));
	// LUT = (~I1&~I2&~I4)|(~ID&I2&~I4)|(I0&I2&I4)|(~I1&~I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4747  */ #(
            .INIT(32'b10001101101011110000010100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4747  (
            .Z (_N10183_178),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_315),
            .I3 (_N10183_576),
            .I4 (_N10183_577));
	// LUT = (I0&I1&I4)|(I0&~I1&~I3)|(~I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4749  (
            .Z (_N10183_180),
            .I0 (_N10183_319_inv),
            .I1 (_N10183_320),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4750  (
            .Z (_N10183_181),
            .I0 (_N10183_322),
            .I1 (_N10183_321),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4751  (
            .Z (_N10183_182),
            .I0 (_N10183_323_inv),
            .I1 (_N10183_324),
            .S (\u_lcd_rgb_char/bcd_data_y [2] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4753  */ #(
            .INIT(32'b11110011111000101101000111000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4753  (
            .Z (_N10183_184),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_328),
            .I3 (_N10183_595),
            .I4 (_N10183_596));
	// LUT = (I0&~I1&I4)|(~I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4754  */ #(
            .INIT(32'b10101010101010100100111101111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4754  (
            .Z (_N10183_185),
            .I0 (_N10183_330),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_1057),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1056));
	// LUT = (~I1&~I3&~I4)|(~I2&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4755  (
            .Z (_N10183_186),
            .I0 (_N10183_331_inv),
            .I1 (_N10183_332),
            .S (\u_lcd_rgb_char/bcd_data_y [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4756  (
            .Z (_N10183_187),
            .I0 (_N10183_333),
            .I1 (_N10183_334),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4757  (
            .Z (_N10183_188),
            .I0 (_N10183_335),
            .I1 (_N10183_336),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4758  */ #(
            .INIT(32'b10110001111101011010000011100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4758  (
            .Z (_N10183_189),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_338),
            .I3 (_N10183_613),
            .I4 (_N10183_614));
	// LUT = (~I0&~I1&I4)|(~I0&I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4759  */ #(
            .INIT(32'b11111100101110000111010000110000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4759  (
            .Z (_N10183_190),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_339),
            .I3 (_N10183_618),
            .I4 (_N10183_619));
	// LUT = (I0&I1&I4)|(~I0&I1&I3)|(~I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4760  (
            .Z (_N10183_191),
            .I0 (_N10183_342),
            .I1 (_N10183_341),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4761  (
            .Z (_N10183_192),
            .I0 (_N10183_343),
            .I1 (_N10183_344),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4762  */ #(
            .INIT(32'b10100000101000110101001101010011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4762  (
            .Z (_N10183_193),
            .I0 (_N10183_629),
            .I1 (_N10183_628),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_630));
	// LUT = (~I1&~I2&~I4)|(~ID&I2&~I4)|(I0&I2&I4)|(~I1&~I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4763  */ #(
            .INIT(32'b10001101101011110000010100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4763  (
            .Z (_N10183_194),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_347),
            .I3 (_N10183_633),
            .I4 (_N10183_634));
	// LUT = (I0&I1&I4)|(I0&~I1&~I3)|(~I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4765  (
            .Z (_N10183_196),
            .I0 (_N10183_350_inv),
            .I1 (_N10183_351),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4766  (
            .Z (_N10183_197),
            .I0 (_N10183_353),
            .I1 (_N10183_352),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4767  (
            .Z (_N10183_198),
            .I0 (_N10183_354_inv),
            .I1 (_N10183_355),
            .S (\u_lcd_rgb_char/bcd_data_x [2] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4769  */ #(
            .INIT(32'b11110011111000101101000111000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4769  (
            .Z (_N10183_200),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_359),
            .I3 (_N10183_651),
            .I4 (_N10183_652));
	// LUT = (I0&~I1&I4)|(~I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4770  */ #(
            .INIT(32'b10101010101010100100111101111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4770  (
            .Z (_N10183_201),
            .I0 (_N10183_361),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_1149),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1148));
	// LUT = (~I1&~I3&~I4)|(~I2&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4771  (
            .Z (_N10183_202),
            .I0 (_N10183_362_inv),
            .I1 (_N10183_363),
            .S (\u_lcd_rgb_char/bcd_data_x [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4772  (
            .Z (_N10183_203),
            .I0 (_N10183_364),
            .I1 (_N10183_365),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4773  (
            .Z (_N10183_204),
            .I0 (_N10183_366),
            .I1 (_N10183_367),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4774  */ #(
            .INIT(32'b10110001111101011010000011100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4774  (
            .Z (_N10183_205),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_369),
            .I3 (_N10183_669),
            .I4 (_N10183_670));
	// LUT = (~I0&~I1&I4)|(~I0&I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4775  */ #(
            .INIT(32'b11111100101110000111010000110000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4775  (
            .Z (_N10183_206),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_370),
            .I3 (_N10183_674),
            .I4 (_N10183_675));
	// LUT = (I0&I1&I4)|(~I0&I1&I3)|(~I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4776  (
            .Z (_N10183_207),
            .I0 (_N10183_373),
            .I1 (_N10183_372),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4777  (
            .Z (_N10183_208),
            .I0 (_N10183_374),
            .I1 (_N10183_375),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4778  */ #(
            .INIT(32'b10100000101000110101001101010011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4778  (
            .Z (_N10183_209),
            .I0 (_N10183_685),
            .I1 (_N10183_684),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_686));
	// LUT = (~I1&~I2&~I4)|(~ID&I2&~I4)|(I0&I2&I4)|(~I1&~I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4779  */ #(
            .INIT(32'b10001101101011110000010100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4779  (
            .Z (_N10183_210),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_378),
            .I3 (_N10183_689),
            .I4 (_N10183_690));
	// LUT = (I0&I1&I4)|(I0&~I1&~I3)|(~I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4781  (
            .Z (_N10183_212),
            .I0 (_N10183_381_inv),
            .I1 (_N10183_382),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4782  (
            .Z (_N10183_213),
            .I0 (_N10183_384),
            .I1 (_N10183_383),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4783  (
            .Z (_N10183_214),
            .I0 (_N10183_385_inv),
            .I1 (_N10183_386),
            .S (\u_lcd_rgb_char/bcd_data_y [6] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4785  */ #(
            .INIT(32'b11110011111000101101000111000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4785  (
            .Z (_N10183_216),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_390),
            .I3 (_N10183_707),
            .I4 (_N10183_708));
	// LUT = (I0&~I1&I4)|(~I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4786  */ #(
            .INIT(32'b10101010101010100100111101111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4786  (
            .Z (_N10183_217),
            .I0 (_N10183_392),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_1240),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1239));
	// LUT = (~I1&~I3&~I4)|(~I2&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4787  (
            .Z (_N10183_218),
            .I0 (_N10183_393_inv),
            .I1 (_N10183_394),
            .S (\u_lcd_rgb_char/bcd_data_y [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4788  (
            .Z (_N10183_219),
            .I0 (_N10183_395),
            .I1 (_N10183_396),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4789  (
            .Z (_N10183_220),
            .I0 (_N10183_397),
            .I1 (_N10183_398),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4790  */ #(
            .INIT(32'b10110001111101011010000011100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4790  (
            .Z (_N10183_221),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_400),
            .I3 (_N10183_725),
            .I4 (_N10183_726));
	// LUT = (~I0&~I1&I4)|(~I0&I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4791  */ #(
            .INIT(32'b11111100101110000111010000110000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4791  (
            .Z (_N10183_222),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_401),
            .I3 (_N10183_730),
            .I4 (_N10183_731));
	// LUT = (I0&I1&I4)|(~I0&I1&I3)|(~I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4792  (
            .Z (_N10183_223),
            .I0 (_N10183_404),
            .I1 (_N10183_403),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4793  (
            .Z (_N10183_224),
            .I0 (_N10183_405),
            .I1 (_N10183_406),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4794  */ #(
            .INIT(32'b10100000101000110101001101010011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4794  (
            .Z (_N10183_225),
            .I0 (_N10183_741),
            .I1 (_N10183_740),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_742));
	// LUT = (~I1&~I2&~I4)|(~ID&I2&~I4)|(I0&I2&I4)|(~I1&~I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4795  */ #(
            .INIT(32'b10001101101011110000010100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4795  (
            .Z (_N10183_226),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_409),
            .I3 (_N10183_745),
            .I4 (_N10183_746));
	// LUT = (I0&I1&I4)|(I0&~I1&~I3)|(~I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4797  (
            .Z (_N10183_228),
            .I0 (_N10183_412_inv),
            .I1 (_N10183_413),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4798  (
            .Z (_N10183_229),
            .I0 (_N10183_415),
            .I1 (_N10183_414),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4799  (
            .Z (_N10183_230),
            .I0 (_N10183_416_inv),
            .I1 (_N10183_417),
            .S (\u_lcd_rgb_char/bcd_data_x [6] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4801  */ #(
            .INIT(32'b11110011111000101101000111000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4801  (
            .Z (_N10183_232),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_421),
            .I3 (_N10183_763),
            .I4 (_N10183_764));
	// LUT = (I0&~I1&I4)|(~I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4802  */ #(
            .INIT(32'b10101010101010100100111101111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4802  (
            .Z (_N10183_233),
            .I0 (_N10183_423),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_1331),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1330));
	// LUT = (~I1&~I3&~I4)|(~I2&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4803  (
            .Z (_N10183_234),
            .I0 (_N10183_424_inv),
            .I1 (_N10183_425),
            .S (\u_lcd_rgb_char/bcd_data_x [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4804  (
            .Z (_N10183_235),
            .I0 (_N10183_426),
            .I1 (_N10183_427),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4805  (
            .Z (_N10183_236),
            .I0 (_N10183_428),
            .I1 (_N10183_429),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4806  */ #(
            .INIT(32'b10110001111101011010000011100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4806  (
            .Z (_N10183_237),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_431),
            .I3 (_N10183_781),
            .I4 (_N10183_782));
	// LUT = (~I0&~I1&I4)|(~I0&I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4807  */ #(
            .INIT(32'b11111100101110000111010000110000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4807  (
            .Z (_N10183_238),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_432),
            .I3 (_N10183_786),
            .I4 (_N10183_787));
	// LUT = (I0&I1&I4)|(~I0&I1&I3)|(~I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4808  (
            .Z (_N10183_239),
            .I0 (_N10183_435),
            .I1 (_N10183_434),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4809  (
            .Z (_N10183_240),
            .I0 (_N10183_436),
            .I1 (_N10183_437),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4810  */ #(
            .INIT(32'b10100000101000110101001101010011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4810  (
            .Z (_N10183_241),
            .I0 (_N10183_797),
            .I1 (_N10183_796),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_798));
	// LUT = (~I1&~I2&~I4)|(~ID&I2&~I4)|(I0&I2&I4)|(~I1&~I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4811  */ #(
            .INIT(32'b10001101101011110000010100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4811  (
            .Z (_N10183_242),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_440),
            .I3 (_N10183_801),
            .I4 (_N10183_802));
	// LUT = (I0&I1&I4)|(I0&~I1&~I3)|(~I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4813  (
            .Z (_N10183_244),
            .I0 (_N10183_443_inv),
            .I1 (_N10183_444),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4814  (
            .Z (_N10183_245),
            .I0 (_N10183_446),
            .I1 (_N10183_445),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4815  (
            .Z (_N10183_246),
            .I0 (_N10183_447_inv),
            .I1 (_N10183_448),
            .S (\u_lcd_rgb_char/bcd_data_y [10] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4817  */ #(
            .INIT(32'b11110011111000101101000111000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4817  (
            .Z (_N10183_248),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_452),
            .I3 (_N10183_819),
            .I4 (_N10183_820));
	// LUT = (I0&~I1&I4)|(~I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4818  */ #(
            .INIT(32'b10101010101010100100111101111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4818  (
            .Z (_N10183_249),
            .I0 (_N10183_454),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_1422),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1421));
	// LUT = (~I1&~I3&~I4)|(~I2&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4819  (
            .Z (_N10183_250),
            .I0 (_N10183_455_inv),
            .I1 (_N10183_456),
            .S (\u_lcd_rgb_char/bcd_data_y [9] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4820  (
            .Z (_N10183_251),
            .I0 (_N10183_457),
            .I1 (_N10183_458),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4821  (
            .Z (_N10183_252),
            .I0 (_N10183_459),
            .I1 (_N10183_460),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4822  */ #(
            .INIT(32'b10110001111101011010000011100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4822  (
            .Z (_N10183_253),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_462),
            .I3 (_N10183_837),
            .I4 (_N10183_838));
	// LUT = (~I0&~I1&I4)|(~I0&I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4823  */ #(
            .INIT(32'b11111100101110000111010000110000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4823  (
            .Z (_N10183_254),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_463),
            .I3 (_N10183_842),
            .I4 (_N10183_843));
	// LUT = (I0&I1&I4)|(~I0&I1&I3)|(~I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4824  (
            .Z (_N10183_255),
            .I0 (_N10183_466),
            .I1 (_N10183_465),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4825  (
            .Z (_N10183_256),
            .I0 (_N10183_467),
            .I1 (_N10183_468),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4826  */ #(
            .INIT(32'b10100000101000110101001101010011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4826  (
            .Z (_N10183_257),
            .I0 (_N10183_853),
            .I1 (_N10183_852),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_854));
	// LUT = (~I1&~I2&~I4)|(~ID&I2&~I4)|(I0&I2&I4)|(~I1&~I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4827  */ #(
            .INIT(32'b10001101101011110000010100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4827  (
            .Z (_N10183_258),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_471),
            .I3 (_N10183_857),
            .I4 (_N10183_858));
	// LUT = (I0&I1&I4)|(I0&~I1&~I3)|(~I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4829  (
            .Z (_N10183_260),
            .I0 (_N10183_474_inv),
            .I1 (_N10183_475),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4830  (
            .Z (_N10183_261),
            .I0 (_N10183_477),
            .I1 (_N10183_476),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4831  (
            .Z (_N10183_262),
            .I0 (_N10183_478_inv),
            .I1 (_N10183_479),
            .S (\u_lcd_rgb_char/bcd_data_x [10] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4833  */ #(
            .INIT(32'b11110011111000101101000111000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4833  (
            .Z (_N10183_264),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_483),
            .I3 (_N10183_875),
            .I4 (_N10183_876));
	// LUT = (I0&~I1&I4)|(~I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4834  */ #(
            .INIT(32'b10101010101010100100111101111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4834  (
            .Z (_N10183_265),
            .I0 (_N10183_485),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_1513),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1512));
	// LUT = (~I1&~I3&~I4)|(~I2&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4835  (
            .Z (_N10183_266),
            .I0 (_N10183_486_inv),
            .I1 (_N10183_487),
            .S (\u_lcd_rgb_char/bcd_data_x [9] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4836  (
            .Z (_N10183_267),
            .I0 (_N10183_488),
            .I1 (_N10183_489),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4837  (
            .Z (_N10183_268),
            .I0 (_N10183_490),
            .I1 (_N10183_491),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4838  */ #(
            .INIT(32'b10110001111101011010000011100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4838  (
            .Z (_N10183_269),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_493),
            .I3 (_N10183_893),
            .I4 (_N10183_894));
	// LUT = (~I0&~I1&I4)|(~I0&I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4839  */ #(
            .INIT(32'b11111100101110000111010000110000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4839  (
            .Z (_N10183_270),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_494),
            .I3 (_N10183_898),
            .I4 (_N10183_899));
	// LUT = (I0&I1&I4)|(~I0&I1&I3)|(~I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4840  (
            .Z (_N10183_271),
            .I0 (_N10183_497),
            .I1 (_N10183_496),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4841  (
            .Z (_N10183_272),
            .I0 (_N10183_498),
            .I1 (_N10183_499),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4842  */ #(
            .INIT(32'b10100000101011110001001100010011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4842  (
            .Z (_N10183_273),
            .I0 (_N10183_909),
            .I1 (_N10183_908),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (_N10183_910),
            .I4 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~I1&~I2&~I4)|(~ID&~I1&~I4)|(~I2&~I3&I4)|(I0&I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4843  */ #(
            .INIT(32'b10001101101011110000010100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4843  (
            .Z (_N10183_274),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_502),
            .I3 (_N10183_913),
            .I4 (_N10183_914));
	// LUT = (I0&I1&I4)|(I0&~I1&~I3)|(~I0&~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4845  (
            .Z (_N10183_276),
            .I0 (_N10183_505_inv),
            .I1 (_N10183_506),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4846  (
            .Z (_N10183_277),
            .I0 (_N10183_508),
            .I1 (_N10183_507),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4847  (
            .Z (_N10183_278),
            .I0 (_N10183_509_inv),
            .I1 (_N10183_510),
            .S (\u_lcd_rgb_char/bcd_data_x [14] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4849  */ #(
            .INIT(32'b11110011111000101101000111000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4849  (
            .Z (_N10183_280),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (_N10183_514),
            .I3 (_N10183_931),
            .I4 (_N10183_932));
	// LUT = (I0&~I1&I4)|(~I0&~I1&I3)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4850  */ #(
            .INIT(32'b10101010101010100100111101111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4850  (
            .Z (_N10183_281),
            .I0 (_N10183_516),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (_N10183_1604),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1603));
	// LUT = (~I1&~I3&~I4)|(~I2&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4851  (
            .Z (_N10183_282),
            .I0 (_N10183_517_inv),
            .I1 (_N10183_518),
            .S (\u_lcd_rgb_char/bcd_data_x [13] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4852  (
            .Z (_N10183_283),
            .I0 (_N10183_519),
            .I1 (_N10183_520),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4853  (
            .Z (_N10183_284),
            .I0 (_N10183_521),
            .I1 (_N10183_522),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4855  */ #(
            .INIT(32'b11111110111011101111111011101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4855  (
            .Z (_N10183_286),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));
	// LUT = (~I2&~I3&~I4)|(I2&I3)|(I1)|(I0) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4857  */ #(
            .INIT(32'b10101010000000110111111101010111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4857  (
            .Z (_N10183_288),
            .I0 (_N10183_953),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));
	// LUT = (~I2&I3&~I4)|(~I1&I3&~I4)|(~ID&~I4)|(I0&I3&I4)|(~I1&~I2&~I3) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_4858_2  */ #(
            .INIT(16'b1111101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4858_2  (
            .Z (_N11860),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (~I3)|(I2)|(~I1)|(I0) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4859  */ #(
            .INIT(32'b11110101000001010100011101000111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4859  (
            .Z (_N10183_290),
            .I0 (_N10183_956),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I3 (_N10183_957),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .ID (_N10183_286));
	// LUT = (~I1&~I2&~I4)|(~ID&I1&~I4)|(I2&I3&I4)|(~I0&~I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4861  */ #(
            .INIT(32'b11000010110000001100000010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4861  (
            .Z (_N10183_292),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I1&~I2&I3&I4)|(I1&I2&I4)|(I1&I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4864_3  */ #(
            .INIT(32'b11111111111111110011011101110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4864_3  (
            .Z (_N10183_295),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I4 (_N10183_962));
	// LUT = (I4)|(~I0&~I3)|(~I0&~I2)|(~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4865  */ #(
            .INIT(32'b11001000110010111111100011111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4865  (
            .Z (_N10183_296),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I3 (_N10183_534),
            .I4 (_N10183_966));
	// LUT = (I2&~I4)|(~I1&~I2&~I3)|(I1&I2)|(I0&I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4869  (
            .Z (_N10183_300),
            .I0 (_N10183_545),
            .I1 (_N10183_546),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4870  */ #(
            .INIT(32'b11001110000000101110111000100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4870  (
            .Z (_N10183_301),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I3 (_N10183_547),
            .I4 (_N10183_1656));
	// LUT = (I0&~I1&~I4)|(I1&I3)|(I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4871  */ #(
            .INIT(32'b11111111111111101111111110101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4871  (
            .Z (_N10183_302),
            .I0 (_N10183_1657),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .ID (_N10183_978));
	// LUT = (ID&~I4)|(I2&I4)|(I1&I4)|(I0&I4)|(I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4875  */ #(
            .INIT(32'b11001111110001011100111111001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4875  (
            .Z (_N10183_306),
            .I0 (_N10183_1673),
            .I1 (_N10183_988),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1674));
	// LUT = (ID&~I2&~I4)|(~I0&~I2&I4)|(~I2&I3)|(I1&I2) ;

    GTP_MUX2LUT8 \u_lcd_rgb_char/u_lcd_display/N9971_4876  (
            .Z (_N10183_307),
            .I0 (_N10183_559),
            .I1 (_N10183_558),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4878  */ #(
            .INIT(32'b11111111101010100101110100001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4878  (
            .Z (_N10183_309),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (_N10183_562),
            .I4 (_N10183_999));
	// LUT = (I0&I4)|(~I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4879  */ #(
            .INIT(32'b11110010101111000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4879  (
            .Z (_N10183_310),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_564));
	// LUT = (~ID&~I4)|(I1&~I2&~I3&I4)|(I2&I3&I4)|(I0&~I1&I3&I4)|(~I1&I2&I4)|(I0&I2&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4880  */ #(
            .INIT(32'b11111101111100111111001110101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4880  (
            .Z (_N10183_311),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .ID (_N10183_1005));
	// LUT = (ID&~I3&~I4)|(~I1&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I2&I3)|(~I0&~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4881_3  */ #(
            .INIT(32'b11111111000011111111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4881_3  (
            .Z (_N10183_312),
            .I0 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_578),
            .I3 (_N10183_1008),
            .I4 (_N10456));
	// LUT = (I0&~I1&~I4)|(I3)|(~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4884  (
            .Z (_N10183_315),
            .I0 (_N10183_574_inv),
            .I1 (_N10183_575),
            .S (\u_lcd_rgb_char/bcd_data_y [1] ));

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_4886  */ #(
            .INIT(8'b11000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4886  (
            .Z (_N10183_317),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&I2)|(~I0&I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4887  (
            .Z (_N10183_318),
            .I0 (_N10183_580),
            .I1 (_N10183_579),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4889  */ #(
            .INIT(32'b11111111001110010010111000101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4889  (
            .Z (_N10183_320),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1031));
	// LUT = (I1&~I2&~I4)|(ID&~I1&~I4)|(I3&I4)|(~I1&I2&I4)|(~I0&~I1&I4)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4890  */ #(
            .INIT(32'b10101010101010101011100011111100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4890  (
            .Z (_N10183_321),
            .I0 (_N10183_586),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_1033),
            .I3 (_N10183_1741),
            .I4 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I1&~I3&~I4)|(~I1&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4891  */ #(
            .INIT(32'b11100100010001000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4891  (
            .Z (_N10183_322),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (_N10183_1037),
            .I2 (_N10183_1748),
            .I3 (_N10183_1749),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_588));
	// LUT = (~ID&~I4)|(I0&I2&I3&I4)|(~I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4893  */ #(
            .INIT(32'b11100111111111111101110111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4893  (
            .Z (_N10183_324),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .ID (_N10183_1044));
	// LUT = (I1&~I4)|(~ID&~I4)|(~I3&I4)|(~I0&~I2&I4)|(I0&~I1&I4)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4894  */ #(
            .INIT(32'b11011101110111011101101111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4894  (
            .Z (_N10183_325),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I3&~I4)|(I0&~I2&~I4)|(~I0&I4)|(~I0&~I1&I3)|(~I0&~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4897  (
            .Z (_N10183_328),
            .I0 (_N10183_597),
            .I1 (_N10183_598),
            .S (\u_lcd_rgb_char/bcd_data_y [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4899  (
            .Z (_N10183_330),
            .I0 (_N10183_601),
            .I1 (_N10183_600),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4901  */ #(
            .INIT(32'b10001101000001011010111100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4901  (
            .Z (_N10183_332),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_605),
            .I3 (_N10183_1066),
            .I4 (_N10183_1067));
	// LUT = (I0&~I1&~I4)|(I0&I1&I3)|(~I0&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4902  */ #(
            .INIT(32'b11111111011111111111111111010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4902  (
            .Z (_N10183_333),
            .I0 (_N10183_2789),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [3] ));
	// LUT = (I1&I2&~I4)|(~I2&I4)|(~I1&I4)|(I3)|(~ID&~I2)|(~I0&I1&I2)|(~ID&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4903  */ #(
            .INIT(32'b11111111110111110010001000000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4903  (
            .Z (_N10183_334),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (_N10183_1803),
            .I4 (_N12282));
	// LUT = (I1&I4)|(~I0&I4)|(I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4904  */ #(
            .INIT(32'b10001000100010000000010001000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4904  (
            .Z (_N10183_335),
            .I0 (_N10183_1076),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (_N10183_1806),
            .I4 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .ID (_N10183_1805));
	// LUT = (~ID&I1&~I3&~I4)|(~ID&I1&~I2&~I4)|(I0&I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4905  */ #(
            .INIT(32'b10101000111111010010000001110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4905  (
            .Z (_N10183_336),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_611),
            .I4 (_N10183_1079));
	// LUT = (I0&I1&I4)|(~I0&~I3)|(I0&~I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4907  */ #(
            .INIT(32'b11001111110001011100111111001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4907  (
            .Z (_N10183_338),
            .I0 (_N10183_1823),
            .I1 (_N10183_1084),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1824));
	// LUT = (ID&~I2&~I4)|(~I0&~I2&I4)|(~I2&I3)|(I1&I2) ;

    GTP_MUX2LUT8 \u_lcd_rgb_char/u_lcd_display/N9971_4908  (
            .Z (_N10183_339),
            .I0 (_N10183_617),
            .I1 (_N10183_616),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4910  */ #(
            .INIT(32'b11111111101010100101110100001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4910  (
            .Z (_N10183_341),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (_N10183_620),
            .I4 (_N10183_1095));
	// LUT = (I0&I4)|(~I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4911  */ #(
            .INIT(32'b11110010101111000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4911  (
            .Z (_N10183_342),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_622));
	// LUT = (~ID&~I4)|(I1&~I2&~I3&I4)|(I2&I3&I4)|(I0&~I1&I3&I4)|(~I1&I2&I4)|(I0&I2&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4912  */ #(
            .INIT(32'b11111101111100111111001110101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4912  (
            .Z (_N10183_343),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .ID (_N10183_1100));
	// LUT = (ID&~I3&~I4)|(~I1&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I2&I3)|(~I0&~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4913_3  */ #(
            .INIT(32'b11111111000011111111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4913_3  (
            .Z (_N10183_344),
            .I0 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_578),
            .I3 (_N10183_1102),
            .I4 (_N10456));
	// LUT = (I0&~I1&~I4)|(I3)|(~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4916  (
            .Z (_N10183_347),
            .I0 (_N10183_631_inv),
            .I1 (_N10183_632),
            .S (\u_lcd_rgb_char/bcd_data_x [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4918  (
            .Z (_N10183_349),
            .I0 (_N10183_636),
            .I1 (_N10183_635),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4920  */ #(
            .INIT(32'b11111111001110010010111000101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4920  (
            .Z (_N10183_351),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N11319_2));
	// LUT = (I1&~I2&~I4)|(ID&~I1&~I4)|(I3&I4)|(~I1&I2&I4)|(~I0&~I1&I4)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4921  */ #(
            .INIT(32'b10101010101010101011100011111100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4921  (
            .Z (_N10183_352),
            .I0 (_N10183_642),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_1126),
            .I3 (_N10183_1886),
            .I4 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I1&~I3&~I4)|(~I1&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4922  */ #(
            .INIT(32'b11100100010001000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4922  (
            .Z (_N10183_353),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (_N10183_1130),
            .I2 (_N10183_1748),
            .I3 (_N10183_1893),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_644));
	// LUT = (~ID&~I4)|(I0&I2&I3&I4)|(~I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4924  */ #(
            .INIT(32'b11100111111111111101110111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4924  (
            .Z (_N10183_355),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .ID (_N10183_1137));
	// LUT = (I1&~I4)|(~ID&~I4)|(~I3&I4)|(~I0&~I2&I4)|(I0&~I1&I4)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4925  */ #(
            .INIT(32'b11011101110111011101101111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4925  (
            .Z (_N10183_356),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I3&~I4)|(I0&~I2&~I4)|(~I0&I4)|(~I0&~I1&I3)|(~I0&~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4928  (
            .Z (_N10183_359),
            .I0 (_N10183_653),
            .I1 (_N10183_654),
            .S (\u_lcd_rgb_char/bcd_data_x [1] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4930  (
            .Z (_N10183_361),
            .I0 (_N10183_657),
            .I1 (_N10183_656),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4932  */ #(
            .INIT(32'b10001101000001011010111100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4932  (
            .Z (_N10183_363),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_661),
            .I3 (_N10183_1157),
            .I4 (_N10183_1158));
	// LUT = (I0&~I1&~I4)|(I0&I1&I3)|(~I0&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4933  */ #(
            .INIT(32'b11111111011111111111111111010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4933  (
            .Z (_N10183_364),
            .I0 (_N10183_2918),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [3] ));
	// LUT = (I1&I2&~I4)|(~I2&I4)|(~I1&I4)|(I3)|(~ID&~I2)|(~I0&I1&I2)|(~ID&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4934  */ #(
            .INIT(32'b11111111110111110010001000000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4934  (
            .Z (_N10183_365),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (_N10183_1803),
            .I4 (_N12284));
	// LUT = (I1&I4)|(~I0&I4)|(I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4935  */ #(
            .INIT(32'b10001000100010000000010001000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4935  (
            .Z (_N10183_366),
            .I0 (_N10183_1167),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_1806),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .ID (_N10183_1943));
	// LUT = (~ID&I1&~I3&~I4)|(~ID&I1&~I2&~I4)|(I0&I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4936  */ #(
            .INIT(32'b10101000111111010010000001110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4936  (
            .Z (_N10183_367),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_667),
            .I4 (_N10183_1170));
	// LUT = (I0&I1&I4)|(~I0&~I3)|(I0&~I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4938  */ #(
            .INIT(32'b11001111110001011100111111001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4938  (
            .Z (_N10183_369),
            .I0 (_N10183_1960),
            .I1 (_N10183_1175),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1961));
	// LUT = (ID&~I2&~I4)|(~I0&~I2&I4)|(~I2&I3)|(I1&I2) ;

    GTP_MUX2LUT8 \u_lcd_rgb_char/u_lcd_display/N9971_4939  (
            .Z (_N10183_370),
            .I0 (_N10183_673),
            .I1 (_N10183_672),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4941  */ #(
            .INIT(32'b11111111101010100101110100001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4941  (
            .Z (_N10183_372),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (_N10183_676),
            .I4 (_N10183_1186));
	// LUT = (I0&I4)|(~I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4942  */ #(
            .INIT(32'b11110010101111000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4942  (
            .Z (_N10183_373),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_678));
	// LUT = (~ID&~I4)|(I1&~I2&~I3&I4)|(I2&I3&I4)|(I0&~I1&I3&I4)|(~I1&I2&I4)|(I0&I2&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4943  */ #(
            .INIT(32'b11111101111100111111001110101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4943  (
            .Z (_N10183_374),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .ID (_N10183_1191));
	// LUT = (ID&~I3&~I4)|(~I1&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I2&I3)|(~I0&~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4944_3  */ #(
            .INIT(32'b11111111000011111111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4944_3  (
            .Z (_N10183_375),
            .I0 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_578),
            .I3 (_N10183_1193),
            .I4 (_N10456));
	// LUT = (I0&~I1&~I4)|(I3)|(~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4947  (
            .Z (_N10183_378),
            .I0 (_N10183_687_inv),
            .I1 (_N10183_688),
            .S (\u_lcd_rgb_char/bcd_data_y [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4949  (
            .Z (_N10183_380),
            .I0 (_N10183_692),
            .I1 (_N10183_691),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4951  */ #(
            .INIT(32'b11111111001110010010111000101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4951  (
            .Z (_N10183_382),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1215));
	// LUT = (I1&~I2&~I4)|(ID&~I1&~I4)|(I3&I4)|(~I1&I2&I4)|(~I0&~I1&I4)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4952  */ #(
            .INIT(32'b10101010101010101011100011111100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4952  (
            .Z (_N10183_383),
            .I0 (_N10183_698),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_1217),
            .I3 (_N10183_2023),
            .I4 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I1&~I3&~I4)|(~I1&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4953  */ #(
            .INIT(32'b11100100010001000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4953  (
            .Z (_N10183_384),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (_N10183_1221),
            .I2 (_N10183_1748),
            .I3 (_N10183_2030),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_700));
	// LUT = (~ID&~I4)|(I0&I2&I3&I4)|(~I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4955  */ #(
            .INIT(32'b11100111111111111101110111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4955  (
            .Z (_N10183_386),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .ID (_N10183_1228));
	// LUT = (I1&~I4)|(~ID&~I4)|(~I3&I4)|(~I0&~I2&I4)|(I0&~I1&I4)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4956  */ #(
            .INIT(32'b11011101110111011101101111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4956  (
            .Z (_N10183_387),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I3&~I4)|(I0&~I2&~I4)|(~I0&I4)|(~I0&~I1&I3)|(~I0&~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4959  (
            .Z (_N10183_390),
            .I0 (_N10183_709),
            .I1 (_N10183_710),
            .S (\u_lcd_rgb_char/bcd_data_y [5] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4961  (
            .Z (_N10183_392),
            .I0 (_N10183_713),
            .I1 (_N10183_712),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4963  */ #(
            .INIT(32'b10001101000001011010111100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4963  (
            .Z (_N10183_394),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_717),
            .I3 (_N10183_1248),
            .I4 (_N10183_1249));
	// LUT = (I0&~I1&~I4)|(I0&I1&I3)|(~I0&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4964  */ #(
            .INIT(32'b11111111011111111111111111010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4964  (
            .Z (_N10183_395),
            .I0 (_N10183_3039),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [7] ));
	// LUT = (I1&I2&~I4)|(~I2&I4)|(~I1&I4)|(I3)|(~ID&~I2)|(~I0&I1&I2)|(~ID&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4965  */ #(
            .INIT(32'b11111111110111110010001000000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4965  (
            .Z (_N10183_396),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (_N10183_1803),
            .I4 (_N12286));
	// LUT = (I1&I4)|(~I0&I4)|(I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4966  */ #(
            .INIT(32'b10001000100010000000010001000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4966  (
            .Z (_N10183_397),
            .I0 (_N10183_1258),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_1806),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .ID (_N10183_2080));
	// LUT = (~ID&I1&~I3&~I4)|(~ID&I1&~I2&~I4)|(I0&I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4967  */ #(
            .INIT(32'b10101000111111010010000001110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4967  (
            .Z (_N10183_398),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_723),
            .I4 (_N10183_1261));
	// LUT = (I0&I1&I4)|(~I0&~I3)|(I0&~I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4969  */ #(
            .INIT(32'b11001111110001011100111111001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4969  (
            .Z (_N10183_400),
            .I0 (_N10183_2097),
            .I1 (_N10183_1266),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_2098));
	// LUT = (ID&~I2&~I4)|(~I0&~I2&I4)|(~I2&I3)|(I1&I2) ;

    GTP_MUX2LUT8 \u_lcd_rgb_char/u_lcd_display/N9971_4970  (
            .Z (_N10183_401),
            .I0 (_N10183_729),
            .I1 (_N10183_728),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4972  */ #(
            .INIT(32'b11111111101010100101110100001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_4972  (
            .Z (_N10183_403),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (_N10183_732),
            .I4 (_N10183_1277));
	// LUT = (I0&I4)|(~I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4973  */ #(
            .INIT(32'b11110010101111000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4973  (
            .Z (_N10183_404),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_734));
	// LUT = (~ID&~I4)|(I1&~I2&~I3&I4)|(I2&I3&I4)|(I0&~I1&I3&I4)|(~I1&I2&I4)|(I0&I2&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4974  */ #(
            .INIT(32'b11111101111100111111001110101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4974  (
            .Z (_N10183_405),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .ID (_N10183_1282));
	// LUT = (ID&~I3&~I4)|(~I1&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I2&I3)|(~I0&~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4975_3  */ #(
            .INIT(32'b11111111000011111111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4975_3  (
            .Z (_N10183_406),
            .I0 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_578),
            .I3 (_N10183_1284),
            .I4 (_N10456));
	// LUT = (I0&~I1&~I4)|(I3)|(~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4978  (
            .Z (_N10183_409),
            .I0 (_N10183_743_inv),
            .I1 (_N10183_744),
            .S (\u_lcd_rgb_char/bcd_data_x [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4980  (
            .Z (_N10183_411),
            .I0 (_N10183_748),
            .I1 (_N10183_747),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4982  */ #(
            .INIT(32'b11111111001110010010111000101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_4982  (
            .Z (_N10183_413),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N11503_2));
	// LUT = (I1&~I2&~I4)|(ID&~I1&~I4)|(I3&I4)|(~I1&I2&I4)|(~I0&~I1&I4)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4983  */ #(
            .INIT(32'b10101010101010101011100011111100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4983  (
            .Z (_N10183_414),
            .I0 (_N10183_754),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_1308),
            .I3 (_N10183_2160),
            .I4 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I1&~I3&~I4)|(~I1&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4984  */ #(
            .INIT(32'b11100100010001000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4984  (
            .Z (_N10183_415),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (_N10183_1312),
            .I2 (_N10183_1748),
            .I3 (_N10183_2167),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_756));
	// LUT = (~ID&~I4)|(I0&I2&I3&I4)|(~I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4986  */ #(
            .INIT(32'b11100111111111111101110111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4986  (
            .Z (_N10183_417),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .ID (_N10183_1319));
	// LUT = (I1&~I4)|(~ID&~I4)|(~I3&I4)|(~I0&~I2&I4)|(I0&~I1&I4)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4987  */ #(
            .INIT(32'b11011101110111011101101111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_4987  (
            .Z (_N10183_418),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I3&~I4)|(I0&~I2&~I4)|(~I0&I4)|(~I0&~I1&I3)|(~I0&~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_4990  (
            .Z (_N10183_421),
            .I0 (_N10183_765),
            .I1 (_N10183_766),
            .S (\u_lcd_rgb_char/bcd_data_x [5] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_4992  (
            .Z (_N10183_423),
            .I0 (_N10183_769),
            .I1 (_N10183_768),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4994  */ #(
            .INIT(32'b10001101000001011010111100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_4994  (
            .Z (_N10183_425),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_773),
            .I3 (_N10183_1339),
            .I4 (_N10183_1340));
	// LUT = (I0&~I1&~I4)|(I0&I1&I3)|(~I0&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4995  */ #(
            .INIT(32'b11111111011111111111111111010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4995  (
            .Z (_N10183_426),
            .I0 (_N10183_3160),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [7] ));
	// LUT = (I1&I2&~I4)|(~I2&I4)|(~I1&I4)|(I3)|(~ID&~I2)|(~I0&I1&I2)|(~ID&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4996  */ #(
            .INIT(32'b11111111110111110010001000000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_4996  (
            .Z (_N10183_427),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (_N10183_1803),
            .I4 (_N12288));
	// LUT = (I1&I4)|(~I0&I4)|(I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_4997  */ #(
            .INIT(32'b10001000100010000000010001000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_4997  (
            .Z (_N10183_428),
            .I0 (_N10183_1349),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_1806),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .ID (_N10183_2217));
	// LUT = (~ID&I1&~I3&~I4)|(~ID&I1&~I2&~I4)|(I0&I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_4998  */ #(
            .INIT(32'b10101000111111010010000001110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_4998  (
            .Z (_N10183_429),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_779),
            .I4 (_N10183_1352));
	// LUT = (I0&I1&I4)|(~I0&~I3)|(I0&~I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5000  */ #(
            .INIT(32'b11001111110001011100111111001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5000  (
            .Z (_N10183_431),
            .I0 (_N10183_2234),
            .I1 (_N10183_1357),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_2235));
	// LUT = (ID&~I2&~I4)|(~I0&~I2&I4)|(~I2&I3)|(I1&I2) ;

    GTP_MUX2LUT8 \u_lcd_rgb_char/u_lcd_display/N9971_5001  (
            .Z (_N10183_432),
            .I0 (_N10183_785),
            .I1 (_N10183_784),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5003  */ #(
            .INIT(32'b11111111101010100101110100001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5003  (
            .Z (_N10183_434),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (_N10183_788),
            .I4 (_N10183_1368));
	// LUT = (I0&I4)|(~I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5004  */ #(
            .INIT(32'b11110010101111000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5004  (
            .Z (_N10183_435),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_790));
	// LUT = (~ID&~I4)|(I1&~I2&~I3&I4)|(I2&I3&I4)|(I0&~I1&I3&I4)|(~I1&I2&I4)|(I0&I2&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5005  */ #(
            .INIT(32'b11111101111100111111001110101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5005  (
            .Z (_N10183_436),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .ID (_N10183_1373));
	// LUT = (ID&~I3&~I4)|(~I1&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I2&I3)|(~I0&~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5006_3  */ #(
            .INIT(32'b11111111000011111111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5006_3  (
            .Z (_N10183_437),
            .I0 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_578),
            .I3 (_N10183_1375),
            .I4 (_N10456));
	// LUT = (I0&~I1&~I4)|(I3)|(~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5009  (
            .Z (_N10183_440),
            .I0 (_N10183_799_inv),
            .I1 (_N10183_800),
            .S (\u_lcd_rgb_char/bcd_data_y [9] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5011  (
            .Z (_N10183_442),
            .I0 (_N10183_804),
            .I1 (_N10183_803),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5013  */ #(
            .INIT(32'b11111111001110010010111000101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5013  (
            .Z (_N10183_444),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1397));
	// LUT = (I1&~I2&~I4)|(ID&~I1&~I4)|(I3&I4)|(~I1&I2&I4)|(~I0&~I1&I4)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5014  */ #(
            .INIT(32'b10101010101010101011100011111100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5014  (
            .Z (_N10183_445),
            .I0 (_N10183_810),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_1399),
            .I3 (_N10183_2297),
            .I4 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I1&~I3&~I4)|(~I1&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5015  */ #(
            .INIT(32'b11100100010001000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5015  (
            .Z (_N10183_446),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (_N10183_1403),
            .I2 (_N10183_1748),
            .I3 (_N10183_2304),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_812));
	// LUT = (~ID&~I4)|(I0&I2&I3&I4)|(~I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5017  */ #(
            .INIT(32'b11100111111111111101110111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5017  (
            .Z (_N10183_448),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .ID (_N10183_1410));
	// LUT = (I1&~I4)|(~ID&~I4)|(~I3&I4)|(~I0&~I2&I4)|(I0&~I1&I4)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5018  */ #(
            .INIT(32'b11011101110111011101101111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5018  (
            .Z (_N10183_449),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I3&~I4)|(I0&~I2&~I4)|(~I0&I4)|(~I0&~I1&I3)|(~I0&~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_5019  */ #(
            .INIT(4'b1011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5019  (
            .Z (_N10183_450),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ));
	// LUT = (~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5021  (
            .Z (_N10183_452),
            .I0 (_N10183_821),
            .I1 (_N10183_822),
            .S (\u_lcd_rgb_char/bcd_data_y [9] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5023  (
            .Z (_N10183_454),
            .I0 (_N10183_825),
            .I1 (_N10183_824),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5025  */ #(
            .INIT(32'b10001101000001011010111100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5025  (
            .Z (_N10183_456),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_829),
            .I3 (_N10183_1430),
            .I4 (_N10183_1431));
	// LUT = (I0&~I1&~I4)|(I0&I1&I3)|(~I0&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5026  */ #(
            .INIT(32'b11111111011111111111111111010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5026  (
            .Z (_N10183_457),
            .I0 (_N10183_3281),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [11] ));
	// LUT = (I1&I2&~I4)|(~I2&I4)|(~I1&I4)|(I3)|(~ID&~I2)|(~I0&I1&I2)|(~ID&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5027  */ #(
            .INIT(32'b11111111110111110010001000000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5027  (
            .Z (_N10183_458),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (_N10183_1803),
            .I4 (_N12290));
	// LUT = (I1&I4)|(~I0&I4)|(I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5028  */ #(
            .INIT(32'b10001000100010000000010001000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5028  (
            .Z (_N10183_459),
            .I0 (_N10183_1440),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_1806),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .ID (_N10183_2354));
	// LUT = (~ID&I1&~I3&~I4)|(~ID&I1&~I2&~I4)|(I0&I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5029  */ #(
            .INIT(32'b10101000111111010010000001110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5029  (
            .Z (_N10183_460),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_835),
            .I4 (_N10183_1443));
	// LUT = (I0&I1&I4)|(~I0&~I3)|(I0&~I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5031  */ #(
            .INIT(32'b11001111110001011100111111001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5031  (
            .Z (_N10183_462),
            .I0 (_N10183_2371),
            .I1 (_N10183_1448),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_2372));
	// LUT = (ID&~I2&~I4)|(~I0&~I2&I4)|(~I2&I3)|(I1&I2) ;

    GTP_MUX2LUT8 \u_lcd_rgb_char/u_lcd_display/N9971_5032  (
            .Z (_N10183_463),
            .I0 (_N10183_841),
            .I1 (_N10183_840),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5034  */ #(
            .INIT(32'b11111111101010100101110100001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5034  (
            .Z (_N10183_465),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (_N10183_844),
            .I4 (_N10183_1459));
	// LUT = (I0&I4)|(~I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5035  */ #(
            .INIT(32'b11110010101111000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5035  (
            .Z (_N10183_466),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_846));
	// LUT = (~ID&~I4)|(I1&~I2&~I3&I4)|(I2&I3&I4)|(I0&~I1&I3&I4)|(~I1&I2&I4)|(I0&I2&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5036  */ #(
            .INIT(32'b11111101111100111111001110101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5036  (
            .Z (_N10183_467),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .ID (_N10183_1464));
	// LUT = (ID&~I3&~I4)|(~I1&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I2&I3)|(~I0&~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5037_3  */ #(
            .INIT(32'b11111111000011111111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5037_3  (
            .Z (_N10183_468),
            .I0 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_578),
            .I3 (_N10183_1466),
            .I4 (_N10456));
	// LUT = (I0&~I1&~I4)|(I3)|(~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5040  (
            .Z (_N10183_471),
            .I0 (_N10183_855_inv),
            .I1 (_N10183_856),
            .S (\u_lcd_rgb_char/bcd_data_x [9] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5042  (
            .Z (_N10183_473),
            .I0 (_N10183_860),
            .I1 (_N10183_859),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5044  */ #(
            .INIT(32'b11111111001110010010111000101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5044  (
            .Z (_N10183_475),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1488));
	// LUT = (I1&~I2&~I4)|(ID&~I1&~I4)|(I3&I4)|(~I1&I2&I4)|(~I0&~I1&I4)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5045  */ #(
            .INIT(32'b10101010101010101011100011111100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5045  (
            .Z (_N10183_476),
            .I0 (_N10183_866),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_1490),
            .I3 (_N10183_2434),
            .I4 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I1&~I3&~I4)|(~I1&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5046  */ #(
            .INIT(32'b11100100010001000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5046  (
            .Z (_N10183_477),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (_N10183_1494),
            .I2 (_N10183_1748),
            .I3 (_N10183_2441),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_868));
	// LUT = (~ID&~I4)|(I0&I2&I3&I4)|(~I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5048  */ #(
            .INIT(32'b11100111111111111101110111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5048  (
            .Z (_N10183_479),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .ID (_N10183_1501));
	// LUT = (I1&~I4)|(~ID&~I4)|(~I3&I4)|(~I0&~I2&I4)|(I0&~I1&I4)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5049  */ #(
            .INIT(32'b11011101110111011101101111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5049  (
            .Z (_N10183_480),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I3&~I4)|(I0&~I2&~I4)|(~I0&I4)|(~I0&~I1&I3)|(~I0&~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_5050  */ #(
            .INIT(4'b1011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5050  (
            .Z (_N10183_481),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ));
	// LUT = (~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5052  (
            .Z (_N10183_483),
            .I0 (_N10183_877),
            .I1 (_N10183_878),
            .S (\u_lcd_rgb_char/bcd_data_x [9] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5054  (
            .Z (_N10183_485),
            .I0 (_N10183_881),
            .I1 (_N10183_880),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5056  */ #(
            .INIT(32'b10001101000001011010111100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5056  (
            .Z (_N10183_487),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_885),
            .I3 (_N10183_1521),
            .I4 (_N10183_1522));
	// LUT = (I0&~I1&~I4)|(I0&I1&I3)|(~I0&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5057  */ #(
            .INIT(32'b11111111011111111111111111010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5057  (
            .Z (_N10183_488),
            .I0 (_N10183_3402),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [11] ));
	// LUT = (I1&I2&~I4)|(~I2&I4)|(~I1&I4)|(I3)|(~ID&~I2)|(~I0&I1&I2)|(~ID&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5058  */ #(
            .INIT(32'b11111111110111110010001000000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5058  (
            .Z (_N10183_489),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (_N10183_1803),
            .I4 (_N12292));
	// LUT = (I1&I4)|(~I0&I4)|(I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5059  */ #(
            .INIT(32'b10001000100010000000010001000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5059  (
            .Z (_N10183_490),
            .I0 (_N10183_1531),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_1806),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .ID (_N10183_2491));
	// LUT = (~ID&I1&~I3&~I4)|(~ID&I1&~I2&~I4)|(I0&I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5060  */ #(
            .INIT(32'b10101000111111010010000001110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5060  (
            .Z (_N10183_491),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_891),
            .I4 (_N10183_1534));
	// LUT = (I0&I1&I4)|(~I0&~I3)|(I0&~I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5062  */ #(
            .INIT(32'b11001111110001011100111111001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5062  (
            .Z (_N10183_493),
            .I0 (_N10183_2508),
            .I1 (_N10183_1539),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_2509));
	// LUT = (ID&~I2&~I4)|(~I0&~I2&I4)|(~I2&I3)|(I1&I2) ;

    GTP_MUX2LUT8 \u_lcd_rgb_char/u_lcd_display/N9971_5063  (
            .Z (_N10183_494),
            .I0 (_N10183_897),
            .I1 (_N10183_896),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5065  */ #(
            .INIT(32'b11111111101010100101110100001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5065  (
            .Z (_N10183_496),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (_N10183_900),
            .I4 (_N10183_1550));
	// LUT = (I0&I4)|(~I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5066  */ #(
            .INIT(32'b11110010101111000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5066  (
            .Z (_N10183_497),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_902));
	// LUT = (~ID&~I4)|(I1&~I2&~I3&I4)|(I2&I3&I4)|(I0&~I1&I3&I4)|(~I1&I2&I4)|(I0&I2&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5067  */ #(
            .INIT(32'b11111101111100111111001110101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5067  (
            .Z (_N10183_498),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .ID (_N10183_1555));
	// LUT = (ID&~I3&~I4)|(~I1&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I2&I3)|(~I0&~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5068_3  */ #(
            .INIT(32'b11111111000011111111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5068_3  (
            .Z (_N10183_499),
            .I0 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_578),
            .I3 (_N10183_1557),
            .I4 (_N10456));
	// LUT = (I0&~I1&~I4)|(I3)|(~I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5071  (
            .Z (_N10183_502),
            .I0 (_N10183_911_inv),
            .I1 (_N10183_912),
            .S (\u_lcd_rgb_char/bcd_data_x [13] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5073  (
            .Z (_N10183_504),
            .I0 (_N10183_916),
            .I1 (_N10183_915),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5075  */ #(
            .INIT(32'b11111111001110010010111000101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5075  (
            .Z (_N10183_506),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1579));
	// LUT = (I1&~I2&~I4)|(ID&~I1&~I4)|(I3&I4)|(~I1&I2&I4)|(~I0&~I1&I4)|(I0&I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5076  */ #(
            .INIT(32'b10101010101010101011100011111100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5076  (
            .Z (_N10183_507),
            .I0 (_N10183_922),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_1581),
            .I3 (_N10183_2571),
            .I4 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I1&~I3&~I4)|(~I1&I2&~I4)|(ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5077  */ #(
            .INIT(32'b11100100010001000101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5077  (
            .Z (_N10183_508),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (_N10183_1585),
            .I2 (_N10183_1748),
            .I3 (_N10183_2578),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_924));
	// LUT = (~ID&~I4)|(I0&I2&I3&I4)|(~I0&I1&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5079  */ #(
            .INIT(32'b11100111111111111101110111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5079  (
            .Z (_N10183_510),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .ID (_N10183_1592));
	// LUT = (I1&~I4)|(~ID&~I4)|(~I3&I4)|(~I0&~I2&I4)|(I0&~I1&I4)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5080  */ #(
            .INIT(32'b11011101110111011101101111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5080  (
            .Z (_N10183_511),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I3&~I4)|(I0&~I2&~I4)|(~I0&I4)|(~I0&~I1&I3)|(~I0&~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_5081  */ #(
            .INIT(4'b1011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5081  (
            .Z (_N10183_512),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ));
	// LUT = (~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5083  (
            .Z (_N10183_514),
            .I0 (_N10183_933),
            .I1 (_N10183_934),
            .S (\u_lcd_rgb_char/bcd_data_x [13] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5085  (
            .Z (_N10183_516),
            .I0 (_N10183_937),
            .I1 (_N10183_936),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5087  */ #(
            .INIT(32'b10001101000001011010111100100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5087  (
            .Z (_N10183_518),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (_N10183_941),
            .I3 (_N10183_1612),
            .I4 (_N10183_1613));
	// LUT = (I0&~I1&~I4)|(I0&I1&I3)|(~I0&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5088  */ #(
            .INIT(32'b11111111011111111111111111010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5088  (
            .Z (_N10183_519),
            .I0 (_N10183_3523),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [15] ));
	// LUT = (I1&I2&~I4)|(~I2&I4)|(~I1&I4)|(I3)|(~ID&~I2)|(~I0&I1&I2)|(~ID&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5089  */ #(
            .INIT(32'b11111111110111110010001000000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5089  (
            .Z (_N10183_520),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (_N10183_1803),
            .I4 (_N12294));
	// LUT = (I1&I4)|(~I0&I4)|(I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5090  */ #(
            .INIT(32'b10001000100010000000010001000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5090  (
            .Z (_N10183_521),
            .I0 (_N10183_1622),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_1806),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .ID (_N10183_2628));
	// LUT = (~ID&I1&~I3&~I4)|(~ID&I1&~I2&~I4)|(I0&I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5091  */ #(
            .INIT(32'b10101000111111010010000001110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5091  (
            .Z (_N10183_522),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_947),
            .I4 (_N10183_1625));
	// LUT = (I0&I1&I4)|(~I0&~I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5096  */ #(
            .INIT(32'b11101010101010101010100011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5096  (
            .Z (_N10183_527),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));
	// LUT = (~I3&~I4)|(I1&I2&I3&I4)|(I0&I4)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5103  */ #(
            .INIT(32'b11111101100111111100111111111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5103  (
            .Z (_N10183_534),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (I2&~I3&~I4)|(~I2&I3&~I4)|(~I2&~I3&I4)|(I2&I3&I4)|(~I0&~I1&~I3)|(I1&I3)|(~I0&~I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5104  */ #(
            .INIT(32'b11111111111111110111011101110001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5104  (
            .Z (_N10183_535),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (_N10183_962));
	// LUT = (I4)|(~I1&I3)|(~I0&I3)|(~I1&I2)|(~I0&I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5111_3  */ #(
            .INIT(32'b10000000000000000000000000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5111_3  (
            .Z (_N10183_542),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = I0&I1&I2&I3&I4 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5112  */ #(
            .INIT(32'b11001101110111001100110011001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5112  (
            .Z (_N10183_543),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (~I0&I2&~I3&I4)|(~I0&~I2&I3&I4)|(I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5113  (
            .Z (_N10183_544),
            .I0 (_N10183_969),
            .I1 (_N10183_970),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5114  */ #(
            .INIT(32'b11110011111100010111000110110001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5114  (
            .Z (_N10183_545),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (~I1&I3&I4)|(I2&I4)|(I0&I2&~I3)|(~I0&I2&I3)|(~I1&I2)|(~I0&~I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5115  */ #(
            .INIT(32'b11111000100100001111000001110000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5115  (
            .Z (_N10183_546),
            .I0 (_N10183_1634),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_1004));
	// LUT = (~I1&I2&~I4)|(~ID&I2&~I4)|(I0&I1&I3&I4)|(I0&I1&I2&I4)|(I2&I3)|(~I0&~I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5116  (
            .Z (_N10183_547),
            .I0 (_N10183_974),
            .I1 (_N10183_975),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5120  */ #(
            .INIT(32'b10000000000000011100000000000011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5120  (
            .Z (_N10183_551),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I1&~I2&~I3&~I4)|(I1&I2&I3&~I4)|(~I0&~I1&~I2&~I3)|(I0&I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5123  (
            .Z (_N10183_554),
            .I0 (_N10183_985_inv),
            .I1 (_N10183_984),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5124  */ #(
            .INIT(32'b11010001110111011110111011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5124  (
            .Z (_N10183_555),
            .I0 (_N11004_2),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .ID (_N10183_1668));
	// LUT = (I1&~I4)|(ID&~I4)|(~I0&~I1&I4)|(I1&~I3)|(I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_5125  */ #(
            .INIT(4'b1101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5125  (
            .Z (_N10183_556),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1)|(~I0) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5127  (
            .Z (_N10183_558),
            .I0 (_N10183_990),
            .I1 (_N10183_991),
            .S (\u_lcd_rgb_char/bcd_data_y [0] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5128  (
            .Z (_N10183_559),
            .I0 (_N10183_993),
            .I1 (_N10183_992),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5130  (
            .Z (_N10183_561),
            .I0 (_N10183_996),
            .I1 (_N10183_995),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5131  */ #(
            .INIT(32'b11110000011111111000111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5131  (
            .Z (_N10183_562),
            .I0 (_N10183_2650),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_556),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(I2&I3&I4)|(~I2&~I3)|(~I1&~I3)|(~I0&~I3)|(ID&I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5133  (
            .Z (_N10183_564),
            .I0 (_N10183_1001_inv),
            .I1 (_N10183_1000),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5140  (
            .Z (_N10183_571),
            .I0 (_N10183_1011_inv),
            .I1 (_N10183_1012),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5141  */ #(
            .INIT(32'b10101111101000111010110010100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5141  (
            .Z (_N10183_572),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_1706),
            .I4 (_N10183_1707));
	// LUT = (~I1&~I2&I4)|(I1&~I2&I3)|(I0&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5142  */ #(
            .INIT(32'b10101010101010101111111101111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5142  (
            .Z (_N10183_573),
            .I0 (_N10183_1015),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [0] ));
	// LUT = (I3&~I4)|(ID&~I2&~I4)|(~ID&I2&~I4)|(ID&~I1&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5144  */ #(
            .INIT(32'b11101110111100111111011111110100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5144  (
            .Z (_N10183_575),
            .I0 (_N12065),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_1716),
            .I3 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~I1&I3&~I4)|(~ID&I1&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&~I3)|(I0&~I1&I3)|(I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5145  (
            .Z (_N10183_576),
            .I0 (_N10183_1020_inv),
            .I1 (_N10183_1021),
            .S (\u_lcd_rgb_char/bcd_data_y [3] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5146  (
            .Z (_N10183_577),
            .I0 (_N10183_1022_inv),
            .I1 (_N10183_1023),
            .S (\u_lcd_rgb_char/bcd_data_y [1] ));

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_5147  */ #(
            .INIT(4'b1101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5147  (
            .Z (_N10183_578),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1)|(~I0) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5148  */ #(
            .INIT(32'b11111110111111001010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5148  (
            .Z (_N10183_579),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .ID (_N10183_1024));
	// LUT = (ID&~I4)|(I0&I3&I4)|(I2&I4)|(I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5149  */ #(
            .INIT(32'b11111111111111111000101000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5149  (
            .Z (_N10183_580),
            .I0 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (_N10183_1026));
	// LUT = (I4)|(I0&~I2&I3)|(I0&I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5155  */ #(
            .INIT(32'b11100100111101011010000010110001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5155  (
            .Z (_N10183_586),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_1036),
            .I3 (_N10183_1742),
            .I4 (_N10183_1743));
	// LUT = (~I0&I1&I4)|(~I0&~I1&~I3)|(I0&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5157  (
            .Z (_N10183_588),
            .I0 (_N10183_1039),
            .I1 (_N10183_1040),
            .S (\u_lcd_rgb_char/bcd_data_y [2] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5158  */ #(
            .INIT(32'b11011111111011100001001100100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5158  (
            .Z (_N10183_589),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_1042));
	// LUT = (I1&I4)|(I0&~I1&~I3)|(~I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5164  (
            .Z (_N10183_595),
            .I0 (_N10183_1049),
            .I1 (_N10183_1048),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5165  (
            .Z (_N10183_596),
            .I0 (_N10183_1051),
            .I1 (_N10183_1050),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5166  */ #(
            .INIT(32'b11111111101101111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5166  (
            .Z (_N10183_597),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1052));
	// LUT = (ID&~I4)|(I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5167_3  */ #(
            .INIT(32'b11111111111110111111111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5167_3  (
            .Z (_N10183_598),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I4)|(I3)|(I2)|(~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5169  (
            .Z (_N10183_600),
            .I0 (_N10183_1058_inv),
            .I1 (_N10183_1059),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5170  (
            .Z (_N10183_601),
            .I0 (_N10183_1061),
            .I1 (_N10183_1060),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5171  (
            .Z (_N10183_602),
            .I0 (_N10183_1062_inv),
            .I1 (_N10183_1063),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5174  */ #(
            .INIT(32'b10101010101010101011111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5174  (
            .Z (_N10183_605),
            .I0 (_N10183_1069),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [2] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(~I1&~I4)|(ID&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5180  (
            .Z (_N10183_611),
            .I0 (_N10183_1078_inv),
            .I1 (_N10183_1077),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5182  (
            .Z (_N10183_613),
            .I0 (_N10183_1081_inv),
            .I1 (_N10183_1080),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5183  */ #(
            .INIT(32'b11010001110111011110111011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5183  (
            .Z (_N10183_614),
            .I0 (_N11190_2),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .ID (_N10183_1818));
	// LUT = (I1&~I4)|(ID&~I4)|(~I0&~I1&I4)|(I1&~I3)|(I1&I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5185  (
            .Z (_N10183_616),
            .I0 (_N10183_1086),
            .I1 (_N10183_1087),
            .S (\u_lcd_rgb_char/bcd_data_x [0] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5186  (
            .Z (_N10183_617),
            .I0 (_N10183_1089),
            .I1 (_N10183_1088),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5188  (
            .Z (_N10183_619),
            .I0 (_N10183_1092),
            .I1 (_N10183_1091),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5189  */ #(
            .INIT(32'b11110000011111111000111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5189  (
            .Z (_N10183_620),
            .I0 (_N10183_2650),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_556),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(I2&I3&I4)|(~I2&~I3)|(~I1&~I3)|(~I0&~I3)|(ID&I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5191  (
            .Z (_N10183_622),
            .I0 (_N10183_1097_inv),
            .I1 (_N10183_1096),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5197  (
            .Z (_N10183_628),
            .I0 (_N10183_1104_inv),
            .I1 (_N10183_1105),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5198  */ #(
            .INIT(32'b10101111101000111010110010100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5198  (
            .Z (_N10183_629),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_1854),
            .I4 (_N10183_1855));
	// LUT = (~I1&~I2&I4)|(I1&~I2&I3)|(I0&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5199  */ #(
            .INIT(32'b10101010101010101111111101111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5199  (
            .Z (_N10183_630),
            .I0 (_N10183_1108),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [0] ));
	// LUT = (I3&~I4)|(ID&~I2&~I4)|(~ID&I2&~I4)|(ID&~I1&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5201  */ #(
            .INIT(32'b11101110111100111111011111110100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5201  (
            .Z (_N10183_632),
            .I0 (_N12065),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_1863),
            .I3 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~I1&I3&~I4)|(~ID&I1&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&~I3)|(I0&~I1&I3)|(I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5202  (
            .Z (_N10183_633),
            .I0 (_N10183_1113_inv),
            .I1 (_N10183_1114),
            .S (\u_lcd_rgb_char/bcd_data_x [3] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5203  (
            .Z (_N10183_634),
            .I0 (_N10183_1115_inv),
            .I1 (_N10183_1116),
            .S (\u_lcd_rgb_char/bcd_data_x [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5204  */ #(
            .INIT(32'b11111110111111001010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5204  (
            .Z (_N10183_635),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .ID (_N10183_1117));
	// LUT = (ID&~I4)|(I0&I3&I4)|(I2&I4)|(I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5205  */ #(
            .INIT(32'b11111111111111111000101000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5205  (
            .Z (_N10183_636),
            .I0 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (_N10183_1119));
	// LUT = (I4)|(I0&~I2&I3)|(I0&I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5211  */ #(
            .INIT(32'b11100100111101011010000010110001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5211  (
            .Z (_N10183_642),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_1129),
            .I3 (_N10183_1887),
            .I4 (_N10183_1888));
	// LUT = (~I0&I1&I4)|(~I0&~I1&~I3)|(I0&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5213  (
            .Z (_N10183_644),
            .I0 (_N10183_1132),
            .I1 (_N10183_1133),
            .S (\u_lcd_rgb_char/bcd_data_x [2] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5214  */ #(
            .INIT(32'b11011111111011100001001100100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5214  (
            .Z (_N10183_645),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_1135));
	// LUT = (I1&I4)|(I0&~I1&~I3)|(~I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5220  (
            .Z (_N10183_651),
            .I0 (_N10183_1142),
            .I1 (_N10183_1141),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5221  (
            .Z (_N10183_652),
            .I0 (_N10183_1144),
            .I1 (_N10183_1143),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5222  */ #(
            .INIT(32'b11111111101101111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5222  (
            .Z (_N10183_653),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1145));
	// LUT = (ID&~I4)|(I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5223_3  */ #(
            .INIT(32'b11111111111110111111111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5223_3  (
            .Z (_N10183_654),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I4)|(I3)|(I2)|(~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5225  (
            .Z (_N10183_656),
            .I0 (_N10183_1150_inv),
            .I1 (_N10183_1151),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5226  (
            .Z (_N10183_657),
            .I0 (_N10183_1153),
            .I1 (_N10183_1152),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5227  (
            .Z (_N10183_658),
            .I0 (_N10183_1154_inv),
            .I1 (_N10183_1155),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5230  */ #(
            .INIT(32'b10101010101010101011111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5230  (
            .Z (_N10183_661),
            .I0 (_N10183_1160),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [2] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(~I1&~I4)|(ID&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5236  (
            .Z (_N10183_667),
            .I0 (_N10183_1169_inv),
            .I1 (_N10183_1168),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5238  (
            .Z (_N10183_669),
            .I0 (_N10183_1172_inv),
            .I1 (_N10183_1171),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5239  */ #(
            .INIT(32'b11010001110111011110111011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5239  (
            .Z (_N10183_670),
            .I0 (_N11502_2),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .ID (_N10183_1955));
	// LUT = (I1&~I4)|(ID&~I4)|(~I0&~I1&I4)|(I1&~I3)|(I1&I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5241  (
            .Z (_N10183_672),
            .I0 (_N10183_1177),
            .I1 (_N10183_1178),
            .S (\u_lcd_rgb_char/bcd_data_y [4] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5242  (
            .Z (_N10183_673),
            .I0 (_N10183_1180),
            .I1 (_N10183_1179),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5244  (
            .Z (_N10183_675),
            .I0 (_N10183_1183),
            .I1 (_N10183_1182),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5245  */ #(
            .INIT(32'b11110000011111111000111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5245  (
            .Z (_N10183_676),
            .I0 (_N10183_2650),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_556),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(I2&I3&I4)|(~I2&~I3)|(~I1&~I3)|(~I0&~I3)|(ID&I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5247  (
            .Z (_N10183_678),
            .I0 (_N10183_1188_inv),
            .I1 (_N10183_1187),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5253  (
            .Z (_N10183_684),
            .I0 (_N10183_1195_inv),
            .I1 (_N10183_1196),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5254  */ #(
            .INIT(32'b10101111101000111010110010100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5254  (
            .Z (_N10183_685),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_1991),
            .I4 (_N10183_1992));
	// LUT = (~I1&~I2&I4)|(I1&~I2&I3)|(I0&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5255  */ #(
            .INIT(32'b10101010101010101111111101111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5255  (
            .Z (_N10183_686),
            .I0 (_N10183_1199),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [4] ));
	// LUT = (I3&~I4)|(ID&~I2&~I4)|(~ID&I2&~I4)|(ID&~I1&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5257  */ #(
            .INIT(32'b11101110111100111111011111110100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5257  (
            .Z (_N10183_688),
            .I0 (_N12065),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_2000),
            .I3 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~I1&I3&~I4)|(~ID&I1&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&~I3)|(I0&~I1&I3)|(I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5258  (
            .Z (_N10183_689),
            .I0 (_N10183_1204_inv),
            .I1 (_N10183_1205),
            .S (\u_lcd_rgb_char/bcd_data_y [7] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5259  (
            .Z (_N10183_690),
            .I0 (_N10183_1206_inv),
            .I1 (_N10183_1207),
            .S (\u_lcd_rgb_char/bcd_data_y [5] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5260  */ #(
            .INIT(32'b11111110111111001010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5260  (
            .Z (_N10183_691),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .ID (_N10183_1208));
	// LUT = (ID&~I4)|(I0&I3&I4)|(I2&I4)|(I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5261  */ #(
            .INIT(32'b11111111111111111000101000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5261  (
            .Z (_N10183_692),
            .I0 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (_N10183_1210));
	// LUT = (I4)|(I0&~I2&I3)|(I0&I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5267  */ #(
            .INIT(32'b11100100111101011010000010110001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5267  (
            .Z (_N10183_698),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_1220),
            .I3 (_N10183_2024),
            .I4 (_N10183_2025));
	// LUT = (~I0&I1&I4)|(~I0&~I1&~I3)|(I0&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5269  (
            .Z (_N10183_700),
            .I0 (_N10183_1223),
            .I1 (_N10183_1224),
            .S (\u_lcd_rgb_char/bcd_data_y [6] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5270  */ #(
            .INIT(32'b11011111111011100001001100100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5270  (
            .Z (_N10183_701),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_1226));
	// LUT = (I1&I4)|(I0&~I1&~I3)|(~I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5276  (
            .Z (_N10183_707),
            .I0 (_N10183_1233),
            .I1 (_N10183_1232),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5277  (
            .Z (_N10183_708),
            .I0 (_N10183_1235),
            .I1 (_N10183_1234),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5278  */ #(
            .INIT(32'b11111111101101111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5278  (
            .Z (_N10183_709),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1236));
	// LUT = (ID&~I4)|(I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5279_3  */ #(
            .INIT(32'b11111111111110111111111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5279_3  (
            .Z (_N10183_710),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I4)|(I3)|(I2)|(~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5281  (
            .Z (_N10183_712),
            .I0 (_N10183_1241_inv),
            .I1 (_N10183_1242),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5282  (
            .Z (_N10183_713),
            .I0 (_N10183_1244),
            .I1 (_N10183_1243),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5283  (
            .Z (_N10183_714),
            .I0 (_N10183_1245_inv),
            .I1 (_N10183_1246),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5286  */ #(
            .INIT(32'b10101010101010101011111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5286  (
            .Z (_N10183_717),
            .I0 (_N10183_1251),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [6] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(~I1&~I4)|(ID&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5292  (
            .Z (_N10183_723),
            .I0 (_N10183_1260_inv),
            .I1 (_N10183_1259),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5294  (
            .Z (_N10183_725),
            .I0 (_N10183_1263_inv),
            .I1 (_N10183_1262),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5295  */ #(
            .INIT(32'b11010001110111011110111011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5295  (
            .Z (_N10183_726),
            .I0 (_N11016_2),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .ID (_N10183_2092));
	// LUT = (I1&~I4)|(ID&~I4)|(~I0&~I1&I4)|(I1&~I3)|(I1&I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5297  (
            .Z (_N10183_728),
            .I0 (_N10183_1268),
            .I1 (_N10183_1269),
            .S (\u_lcd_rgb_char/bcd_data_x [4] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5298  (
            .Z (_N10183_729),
            .I0 (_N10183_1271),
            .I1 (_N10183_1270),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5300  (
            .Z (_N10183_731),
            .I0 (_N10183_1274),
            .I1 (_N10183_1273),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5301  */ #(
            .INIT(32'b11110000011111111000111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5301  (
            .Z (_N10183_732),
            .I0 (_N10183_2650),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_556),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(I2&I3&I4)|(~I2&~I3)|(~I1&~I3)|(~I0&~I3)|(ID&I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5303  (
            .Z (_N10183_734),
            .I0 (_N10183_1279_inv),
            .I1 (_N10183_1278),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5309  (
            .Z (_N10183_740),
            .I0 (_N10183_1286_inv),
            .I1 (_N10183_1287),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5310  */ #(
            .INIT(32'b10101111101000111010110010100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5310  (
            .Z (_N10183_741),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_2128),
            .I4 (_N10183_2129));
	// LUT = (~I1&~I2&I4)|(I1&~I2&I3)|(I0&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5311  */ #(
            .INIT(32'b10101010101010101111111101111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5311  (
            .Z (_N10183_742),
            .I0 (_N10183_1290),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [4] ));
	// LUT = (I3&~I4)|(ID&~I2&~I4)|(~ID&I2&~I4)|(ID&~I1&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5313  */ #(
            .INIT(32'b11101110111100111111011111110100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5313  (
            .Z (_N10183_744),
            .I0 (_N12065),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_2137),
            .I3 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~I1&I3&~I4)|(~ID&I1&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&~I3)|(I0&~I1&I3)|(I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5314  (
            .Z (_N10183_745),
            .I0 (_N10183_1295_inv),
            .I1 (_N10183_1296),
            .S (\u_lcd_rgb_char/bcd_data_x [7] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5315  (
            .Z (_N10183_746),
            .I0 (_N10183_1297_inv),
            .I1 (_N10183_1298),
            .S (\u_lcd_rgb_char/bcd_data_x [5] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5316  */ #(
            .INIT(32'b11111110111111001010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5316  (
            .Z (_N10183_747),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .ID (_N10183_1299));
	// LUT = (ID&~I4)|(I0&I3&I4)|(I2&I4)|(I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5317  */ #(
            .INIT(32'b11111111111111111000101000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5317  (
            .Z (_N10183_748),
            .I0 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (_N10183_1301));
	// LUT = (I4)|(I0&~I2&I3)|(I0&I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5323  */ #(
            .INIT(32'b11100100111101011010000010110001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5323  (
            .Z (_N10183_754),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_1311),
            .I3 (_N10183_2161),
            .I4 (_N10183_2162));
	// LUT = (~I0&I1&I4)|(~I0&~I1&~I3)|(I0&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5325  (
            .Z (_N10183_756),
            .I0 (_N10183_1314),
            .I1 (_N10183_1315),
            .S (\u_lcd_rgb_char/bcd_data_x [6] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5326  */ #(
            .INIT(32'b11011111111011100001001100100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5326  (
            .Z (_N10183_757),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_1317));
	// LUT = (I1&I4)|(I0&~I1&~I3)|(~I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5332  (
            .Z (_N10183_763),
            .I0 (_N10183_1324),
            .I1 (_N10183_1323),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5333  (
            .Z (_N10183_764),
            .I0 (_N10183_1326),
            .I1 (_N10183_1325),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5334  */ #(
            .INIT(32'b11111111101101111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5334  (
            .Z (_N10183_765),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1327));
	// LUT = (ID&~I4)|(I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5335_3  */ #(
            .INIT(32'b11111111111110111111111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5335_3  (
            .Z (_N10183_766),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I4)|(I3)|(I2)|(~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5337  (
            .Z (_N10183_768),
            .I0 (_N10183_1332_inv),
            .I1 (_N10183_1333),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5338  (
            .Z (_N10183_769),
            .I0 (_N10183_1335),
            .I1 (_N10183_1334),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5339  (
            .Z (_N10183_770),
            .I0 (_N10183_1336_inv),
            .I1 (_N10183_1337),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5342  */ #(
            .INIT(32'b10101010101010101011111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5342  (
            .Z (_N10183_773),
            .I0 (_N10183_1342),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [6] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(~I1&~I4)|(ID&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5348  (
            .Z (_N10183_779),
            .I0 (_N10183_1351_inv),
            .I1 (_N10183_1350),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5350  (
            .Z (_N10183_781),
            .I0 (_N10183_1354_inv),
            .I1 (_N10183_1353),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5351  */ #(
            .INIT(32'b11010001110111011110111011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5351  (
            .Z (_N10183_782),
            .I0 (_N11168_2),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .ID (_N10183_2229));
	// LUT = (I1&~I4)|(ID&~I4)|(~I0&~I1&I4)|(I1&~I3)|(I1&I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5353  (
            .Z (_N10183_784),
            .I0 (_N10183_1359),
            .I1 (_N10183_1360),
            .S (\u_lcd_rgb_char/bcd_data_y [8] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5354  (
            .Z (_N10183_785),
            .I0 (_N10183_1362),
            .I1 (_N10183_1361),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5356  (
            .Z (_N10183_787),
            .I0 (_N10183_1365),
            .I1 (_N10183_1364),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5357  */ #(
            .INIT(32'b11110000011111111000111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5357  (
            .Z (_N10183_788),
            .I0 (_N10183_2650),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_556),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(I2&I3&I4)|(~I2&~I3)|(~I1&~I3)|(~I0&~I3)|(ID&I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5359  (
            .Z (_N10183_790),
            .I0 (_N10183_1370_inv),
            .I1 (_N10183_1369),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5365  (
            .Z (_N10183_796),
            .I0 (_N10183_1377_inv),
            .I1 (_N10183_1378),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5366  */ #(
            .INIT(32'b10101111101000111010110010100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5366  (
            .Z (_N10183_797),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_2265),
            .I4 (_N10183_2266));
	// LUT = (~I1&~I2&I4)|(I1&~I2&I3)|(I0&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5367  */ #(
            .INIT(32'b10101010101010101111111101111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5367  (
            .Z (_N10183_798),
            .I0 (_N10183_1381),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [8] ));
	// LUT = (I3&~I4)|(ID&~I2&~I4)|(~ID&I2&~I4)|(ID&~I1&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5369  */ #(
            .INIT(32'b11101110111100111111011111110100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5369  (
            .Z (_N10183_800),
            .I0 (_N12065),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_2274),
            .I3 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~I1&I3&~I4)|(~ID&I1&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&~I3)|(I0&~I1&I3)|(I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5370  (
            .Z (_N10183_801),
            .I0 (_N10183_1386_inv),
            .I1 (_N10183_1387),
            .S (\u_lcd_rgb_char/bcd_data_y [11] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5371  (
            .Z (_N10183_802),
            .I0 (_N10183_1388_inv),
            .I1 (_N10183_1389),
            .S (\u_lcd_rgb_char/bcd_data_y [9] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5372  */ #(
            .INIT(32'b11111110111111001010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5372  (
            .Z (_N10183_803),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .ID (_N10183_1390));
	// LUT = (ID&~I4)|(I0&I3&I4)|(I2&I4)|(I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5373  */ #(
            .INIT(32'b11111111111111111000101000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5373  (
            .Z (_N10183_804),
            .I0 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (_N10183_1392));
	// LUT = (I4)|(I0&~I2&I3)|(I0&I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5379  */ #(
            .INIT(32'b11100100111101011010000010110001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5379  (
            .Z (_N10183_810),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_1402),
            .I3 (_N10183_2298),
            .I4 (_N10183_2299));
	// LUT = (~I0&I1&I4)|(~I0&~I1&~I3)|(I0&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5381  (
            .Z (_N10183_812),
            .I0 (_N10183_1405),
            .I1 (_N10183_1406),
            .S (\u_lcd_rgb_char/bcd_data_y [10] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5382  */ #(
            .INIT(32'b11011111111011100001001100100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5382  (
            .Z (_N10183_813),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_1408));
	// LUT = (I1&I4)|(I0&~I1&~I3)|(~I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5388  (
            .Z (_N10183_819),
            .I0 (_N10183_1415),
            .I1 (_N10183_1414),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5389  (
            .Z (_N10183_820),
            .I0 (_N10183_1417),
            .I1 (_N10183_1416),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5390  */ #(
            .INIT(32'b11111111101101111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5390  (
            .Z (_N10183_821),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1418));
	// LUT = (ID&~I4)|(I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5391_3  */ #(
            .INIT(32'b11111111111110111111111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5391_3  (
            .Z (_N10183_822),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I4)|(I3)|(I2)|(~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5393  (
            .Z (_N10183_824),
            .I0 (_N10183_1423_inv),
            .I1 (_N10183_1424),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5394  (
            .Z (_N10183_825),
            .I0 (_N10183_1426),
            .I1 (_N10183_1425),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5395  (
            .Z (_N10183_826),
            .I0 (_N10183_1427_inv),
            .I1 (_N10183_1428),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5398  */ #(
            .INIT(32'b10101010101010101011111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5398  (
            .Z (_N10183_829),
            .I0 (_N10183_1433),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [10] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(~I1&~I4)|(ID&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5404  (
            .Z (_N10183_835),
            .I0 (_N10183_1442_inv),
            .I1 (_N10183_1441),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5406  (
            .Z (_N10183_837),
            .I0 (_N10183_1445_inv),
            .I1 (_N10183_1444),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5407  */ #(
            .INIT(32'b11010001110111011110111011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5407  (
            .Z (_N10183_838),
            .I0 (_N11489_2),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .ID (_N10183_2366));
	// LUT = (I1&~I4)|(ID&~I4)|(~I0&~I1&I4)|(I1&~I3)|(I1&I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5409  (
            .Z (_N10183_840),
            .I0 (_N10183_1450),
            .I1 (_N10183_1451),
            .S (\u_lcd_rgb_char/bcd_data_x [8] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5410  (
            .Z (_N10183_841),
            .I0 (_N10183_1453),
            .I1 (_N10183_1452),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5412  (
            .Z (_N10183_843),
            .I0 (_N10183_1456),
            .I1 (_N10183_1455),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5413  */ #(
            .INIT(32'b11110000011111111000111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5413  (
            .Z (_N10183_844),
            .I0 (_N10183_2650),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_556),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(I2&I3&I4)|(~I2&~I3)|(~I1&~I3)|(~I0&~I3)|(ID&I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5415  (
            .Z (_N10183_846),
            .I0 (_N10183_1461_inv),
            .I1 (_N10183_1460),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5421  (
            .Z (_N10183_852),
            .I0 (_N10183_1468_inv),
            .I1 (_N10183_1469),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5422  */ #(
            .INIT(32'b10101111101000111010110010100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5422  (
            .Z (_N10183_853),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (_N10183_2402),
            .I4 (_N10183_2403));
	// LUT = (~I1&~I2&I4)|(I1&~I2&I3)|(I0&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5423  */ #(
            .INIT(32'b10101010101010101111111101111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5423  (
            .Z (_N10183_854),
            .I0 (_N10183_1472),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [8] ));
	// LUT = (I3&~I4)|(ID&~I2&~I4)|(~ID&I2&~I4)|(ID&~I1&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5425  */ #(
            .INIT(32'b11101110111100111111011111110100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5425  (
            .Z (_N10183_856),
            .I0 (_N12065),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_2411),
            .I3 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~I1&I3&~I4)|(~ID&I1&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&~I3)|(I0&~I1&I3)|(I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5426  (
            .Z (_N10183_857),
            .I0 (_N10183_1477_inv),
            .I1 (_N10183_1478),
            .S (\u_lcd_rgb_char/bcd_data_x [11] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5427  (
            .Z (_N10183_858),
            .I0 (_N10183_1479_inv),
            .I1 (_N10183_1480),
            .S (\u_lcd_rgb_char/bcd_data_x [9] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5428  */ #(
            .INIT(32'b11111110111111001010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5428  (
            .Z (_N10183_859),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .ID (_N10183_1481));
	// LUT = (ID&~I4)|(I0&I3&I4)|(I2&I4)|(I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5429  */ #(
            .INIT(32'b11111111111111111000101000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5429  (
            .Z (_N10183_860),
            .I0 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (_N10183_1483));
	// LUT = (I4)|(I0&~I2&I3)|(I0&I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5435  */ #(
            .INIT(32'b11100100111101011010000010110001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5435  (
            .Z (_N10183_866),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_1493),
            .I3 (_N10183_2435),
            .I4 (_N10183_2436));
	// LUT = (~I0&I1&I4)|(~I0&~I1&~I3)|(I0&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5437  (
            .Z (_N10183_868),
            .I0 (_N10183_1496),
            .I1 (_N10183_1497),
            .S (\u_lcd_rgb_char/bcd_data_x [10] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5438  */ #(
            .INIT(32'b11011111111011100001001100100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5438  (
            .Z (_N10183_869),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_1499));
	// LUT = (I1&I4)|(I0&~I1&~I3)|(~I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5444  (
            .Z (_N10183_875),
            .I0 (_N10183_1506),
            .I1 (_N10183_1505),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5445  (
            .Z (_N10183_876),
            .I0 (_N10183_1508),
            .I1 (_N10183_1507),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5446  */ #(
            .INIT(32'b11111111101101111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5446  (
            .Z (_N10183_877),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1509));
	// LUT = (ID&~I4)|(I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5447_3  */ #(
            .INIT(32'b11111111111110111111111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5447_3  (
            .Z (_N10183_878),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I4)|(I3)|(I2)|(~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5449  (
            .Z (_N10183_880),
            .I0 (_N10183_1514_inv),
            .I1 (_N10183_1515),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5450  (
            .Z (_N10183_881),
            .I0 (_N10183_1517),
            .I1 (_N10183_1516),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5451  (
            .Z (_N10183_882),
            .I0 (_N10183_1518_inv),
            .I1 (_N10183_1519),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5454  */ #(
            .INIT(32'b10101010101010101011111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5454  (
            .Z (_N10183_885),
            .I0 (_N10183_1524),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [10] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(~I1&~I4)|(ID&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5460  (
            .Z (_N10183_891),
            .I0 (_N10183_1533_inv),
            .I1 (_N10183_1532),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5462  (
            .Z (_N10183_893),
            .I0 (_N10183_1536_inv),
            .I1 (_N10183_1535),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5463  */ #(
            .INIT(32'b11010001110111011110111011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5463  (
            .Z (_N10183_894),
            .I0 (_N11179_2),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .ID (_N10183_2503));
	// LUT = (I1&~I4)|(ID&~I4)|(~I0&~I1&I4)|(I1&~I3)|(I1&I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5465  (
            .Z (_N10183_896),
            .I0 (_N10183_1541),
            .I1 (_N10183_1542),
            .S (\u_lcd_rgb_char/bcd_data_x [12] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5466  (
            .Z (_N10183_897),
            .I0 (_N10183_1544),
            .I1 (_N10183_1543),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5468  (
            .Z (_N10183_899),
            .I0 (_N10183_1547),
            .I1 (_N10183_1546),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5469  */ #(
            .INIT(32'b11110000011111111000111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5469  (
            .Z (_N10183_900),
            .I0 (_N10183_2650),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_556),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .ID (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(I2&I3&I4)|(~I2&~I3)|(~I1&~I3)|(~I0&~I3)|(ID&I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5471  (
            .Z (_N10183_902),
            .I0 (_N10183_1552_inv),
            .I1 (_N10183_1551),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5477  (
            .Z (_N10183_908),
            .I0 (_N10183_1559_inv),
            .I1 (_N10183_1560),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_5478  */ #(
            .INIT(8'b10111000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5478  (
            .Z (_N10183_909),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (_N10183_1561));
	// LUT = (~I1&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5479  */ #(
            .INIT(32'b10101010101010101111111101111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5479  (
            .Z (_N10183_910),
            .I0 (_N10183_1563),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [12] ));
	// LUT = (I3&~I4)|(ID&~I2&~I4)|(~ID&I2&~I4)|(ID&~I1&~I4)|(~ID&I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5481  */ #(
            .INIT(32'b11101110111100111111011111110100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5481  (
            .Z (_N10183_912),
            .I0 (_N12065),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (_N10183_2548),
            .I3 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (~I1&I3&~I4)|(~ID&I1&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&~I3)|(I0&~I1&I3)|(I1&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5482  (
            .Z (_N10183_913),
            .I0 (_N10183_1568_inv),
            .I1 (_N10183_1569),
            .S (\u_lcd_rgb_char/bcd_data_x [15] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5483  (
            .Z (_N10183_914),
            .I0 (_N10183_1570_inv),
            .I1 (_N10183_1571),
            .S (\u_lcd_rgb_char/bcd_data_x [13] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5484  */ #(
            .INIT(32'b11111110111111001010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5484  (
            .Z (_N10183_915),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .ID (_N10183_1572));
	// LUT = (ID&~I4)|(I0&I3&I4)|(I2&I4)|(I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5485  */ #(
            .INIT(32'b11111111111111111000101000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5485  (
            .Z (_N10183_916),
            .I0 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (_N10183_1574));
	// LUT = (I4)|(I0&~I2&I3)|(I0&I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5491  */ #(
            .INIT(32'b11100100111101011010000010110001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5491  (
            .Z (_N10183_922),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I2 (_N10183_1584),
            .I3 (_N10183_2572),
            .I4 (_N10183_2573));
	// LUT = (~I0&I1&I4)|(~I0&~I1&~I3)|(I0&I2) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5493  (
            .Z (_N10183_924),
            .I0 (_N10183_1587),
            .I1 (_N10183_1588),
            .S (\u_lcd_rgb_char/bcd_data_x [14] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5494  */ #(
            .INIT(32'b11011111111011100001001100100010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5494  (
            .Z (_N10183_925),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (_N10183_1590));
	// LUT = (I1&I4)|(I0&~I1&~I3)|(~I0&~I1&I3)|(I0&~I1&~I2) ;

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5500  (
            .Z (_N10183_931),
            .I0 (_N10183_1597),
            .I1 (_N10183_1596),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT7 \u_lcd_rgb_char/u_lcd_display/N9971_5501  (
            .Z (_N10183_932),
            .I0 (_N10183_1599),
            .I1 (_N10183_1598),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5502  */ #(
            .INIT(32'b11111111101101111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5502  (
            .Z (_N10183_933),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1600));
	// LUT = (ID&~I4)|(I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5503_3  */ #(
            .INIT(32'b11111111111110111111111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5503_3  (
            .Z (_N10183_934),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I4)|(I3)|(I2)|(~I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5505  (
            .Z (_N10183_936),
            .I0 (_N10183_1605_inv),
            .I1 (_N10183_1606),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5506  (
            .Z (_N10183_937),
            .I0 (_N10183_1608),
            .I1 (_N10183_1607),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5507  (
            .Z (_N10183_938),
            .I0 (_N10183_1609_inv),
            .I1 (_N10183_1610),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5510  */ #(
            .INIT(32'b10101010101010101011111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5510  (
            .Z (_N10183_941),
            .I0 (_N10183_1615),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [14] ));
	// LUT = (~I3&~I4)|(~I2&~I4)|(~I1&~I4)|(ID&~I4)|(I0&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5516  (
            .Z (_N10183_947),
            .I0 (_N10183_1624_inv),
            .I1 (_N10183_1623),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5522  */ #(
            .INIT(32'b10111011101110110111111111110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5522  (
            .Z (_N10183_953),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ));
	// LUT = (~I0&~I4)|(I0&I4)|(I0&I2&~I3)|(I0&~I2&I3)|(~I1&I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5526  */ #(
            .INIT(32'b11111111101110111011101100110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5526  (
            .Z (_N10183_957),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (~I0&~I2&~I3&~I4)|(I3&I4)|(I0&I4)|(I0&I3)|(~I1) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_5531  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5531  (
            .Z (_N10183_962),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [6] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5533  */ #(
            .INIT(32'b11111110111011101100111110001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5533  (
            .Z (_N10183_964),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I2&I3&~I4)|(I2&I3&I4)|(I1&I4)|(I0&I4)|(I1&I3)|(I1&~I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5535  */ #(
            .INIT(32'b10001000100001000100001000100001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5535  (
            .Z (_N10183_966),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (~I0&~I1&~I2&~I3&~I4)|(I0&~I1&I2&~I3&~I4)|(I0&~I1&~I2&I3&~I4)|(~I0&I1&I2&I3&~I4)|(~I0&I1&~I2&~I3&I4)|(I0&I1&I3&I4)|(I0&I1&I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5538  */ #(
            .INIT(32'b11111111111111111111111111110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5538  (
            .Z (_N10183_969),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (I4)|(I3)|(I2)|(~I1)|(~I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5539  */ #(
            .INIT(32'b10101110110011001100110111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5539  (
            .Z (_N10183_970),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (~I2&~I3&~I4)|(~I0&~I3&~I4)|(~I0&~I2&~I4)|(I1&~I4)|(I0&I3&I4)|(I1&~I3)|(I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5543_3  */ #(
            .INIT(32'b11111111111111111101110111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5543_3  (
            .Z (_N10183_974),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (I4)|(~I2&~I3)|(I1)|(~I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5544_3  */ #(
            .INIT(32'b11101100110111011111111111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5544_3  (
            .Z (_N10183_975),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (~I4)|(~I0&~I3)|(I0&I2&I3)|(I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5547  */ #(
            .INIT(32'b11001101110110001000000000000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5547  (
            .Z (_N10183_978),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I0&I2&~I3&I4)|(~I0&~I2&I3&I4)|(I1&I2&I4)|(I0&I1&I4)|(I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5552  */ #(
            .INIT(32'b10000011110000011110111111100111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5552  (
            .Z (_N10183_983),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I0&I3&~I4)|(I0&~I1&~I4)|(~I0&I1&~I4)|(I1&I2&~I3)|(~I1&~I2&I3)|(~I0&~I1&~I2)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5553  */ #(
            .INIT(32'b10111011000000010010000110111010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5553  (
            .Z (_N10183_984),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&I2&~I3&~I4)|(I0&~I3&~I4)|(~I1&I3&I4)|(I0&I3&I4)|(~I0&~I1&~I2&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5557  (
            .Z (_N10183_988),
            .I0 (_N10183_1672),
            .I1 (_N10183_1671),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5559  (
            .Z (_N10183_990),
            .I0 (_N10183_1675),
            .I1 (_N10183_1676),
            .S (\u_lcd_rgb_char/bcd_data_y [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5560  (
            .Z (_N10183_991),
            .I0 (_N10183_1677),
            .I1 (_N10183_1678),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5561  (
            .Z (_N10183_992),
            .I0 (_N10183_1680),
            .I1 (_N10183_1679),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5562  (
            .Z (_N10183_993),
            .I0 (_N10183_1682),
            .I1 (_N10183_1681),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5564  */ #(
            .INIT(32'b11111110111110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5564  (
            .Z (_N10183_995),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1685));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5565  */ #(
            .INIT(32'b11101111111111111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5565  (
            .Z (_N10183_996),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .ID (_N10183_1686));
	// LUT = (ID&~I4)|(~I3&I4)|(~I2&I4)|(I1&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5568  */ #(
            .INIT(32'b10111111110110011101101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5568  (
            .Z (_N10183_999),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&I2&~I4)|(~I2&I3&I4)|(I0&I3&I4)|(~I0&I2&~I3)|(I0&~I2&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5569  */ #(
            .INIT(32'b10011000010110100111010011000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5569  (
            .Z (_N10183_1000),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&I2&~I3&~I4)|(~I1&I2&I3&~I4)|(~I0&I1&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(~I0&I1&I2&~I3) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_5573  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5573  (
            .Z (_N10183_1004),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5574  */ #(
            .INIT(32'b10111011111100111011101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5574  (
            .Z (_N10183_1005),
            .I0 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(I2&~I3)|(I0&I3)|(~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5577  */ #(
            .INIT(32'b10011111100111101111100111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5577  (
            .Z (_N10183_1008),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2&~I4)|(I1&~I2&I4)|(I0&~I2&I4)|(I1&~I2&~I3)|(I0&~I2&~I3)|(~I0&~I1&I3)|(~I0&~I1&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5581  */ #(
            .INIT(32'b11101000111111101110111111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5581  (
            .Z (_N10183_1012),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (_N10183_2710));
	// LUT = (~I2&~I4)|(ID&~I4)|(I2&~I3&I4)|(I0&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5584  */ #(
            .INIT(32'b11101100111011001101101110011011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5584  (
            .Z (_N10183_1015),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I2&~I4)|(~I0&~I1&~I4)|(I0&I2&I4)|(I1&I4)|(I1&I2&I3)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5590  */ #(
            .INIT(32'b11110111110001111101001111110011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5590  (
            .Z (_N10183_1021),
            .I0 (_N10183_2712),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .ID (_N10183_2642));
	// LUT = (~I1&~I3&~I4)|(~I1&I3&I4)|(~I0&I1&I4)|(~ID&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5592  */ #(
            .INIT(32'b11001100001100110000110100100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5592  (
            .Z (_N10183_1023),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I2&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I0&~I1&I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5593  */ #(
            .INIT(32'b11110110111111101111100010011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5593  (
            .Z (_N10183_1024),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I4)|(I0&~I1&I4)|(~I0&I1&I4)|(I0&I1&~I3)|(I2&I3)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5595  */ #(
            .INIT(32'b11101111011011110000100101101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5595  (
            .Z (_N10183_1026),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I0&I1&I4)|(I0&~I1&~I3)|(~I0&I1&~I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5597  */ #(
            .INIT(32'b10100101101001010001000100000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5597  (
            .Z (_N10183_1028),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I3&~I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5598_3  */ #(
            .INIT(32'b11001100000100011111111111111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5598_3  (
            .Z (_N10183_1029),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1004));
	// LUT = (I3&~I4)|(I2&~I4)|(I1&~I4)|(~ID&~I4)|(~I0&~I1&~I3&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5599  */ #(
            .INIT(32'b11110101000100010100010011110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5599  (
            .Z (_N10183_1030),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I2&~I3&~I4)|(~I0&I1&~I4)|(I2&I3&I4)|(~I0&~I1&I4)|(~I0&~I1&~I3)|(~I0&I1&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5602  (
            .Z (_N10183_1033),
            .I0 (_N10183_1739),
            .I1 (_N10183_1740),
            .S (\u_lcd_rgb_char/bcd_data_y [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5605  */ #(
            .INIT(32'b11111111101100110101100111101101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5605  (
            .Z (_N10183_1036),
            .I0 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(ID&~I1&I2&~I3)|(I0&ID&I2&~I3)|(ID&I1&~I2&I3)|(~ID&I2&I3)|(~ID&~I1&~I2)|(I0&~ID&I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5606  */ #(
            .INIT(32'b10101010101010101100111011001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5606  (
            .Z (_N10183_1037),
            .I0 (_N10183_1747),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [1] ));
	// LUT = (ID&~I2&I3&~I4)|(I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5608  */ #(
            .INIT(32'b11011110000100101101110000010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5608  (
            .Z (_N10183_1039),
            .I0 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I3 (_N10183_1750),
            .I4 (_N10183_1748),
            .ID (\u_lcd_rgb_char/bcd_data_y [0] ));
	// LUT = (~ID&~I1&I2&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5609  */ #(
            .INIT(32'b10101000011010000000001000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5609  (
            .Z (_N10183_1040),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&I1&I2&~I3&I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(I0&~I1&I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5611  */ #(
            .INIT(32'b10100101111100011110001001011010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5611  (
            .Z (_N10183_1042),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I3&~I4)|(I0&~I1&~I2&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&I2&I4)|(~I0&I2&~I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5612  */ #(
            .INIT(32'b11101010110010001100101010010100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5612  (
            .Z (_N10183_1043),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I0&I3&I4)|(I1&I2&I4)|(I0&I1&I4)|(I0&~I2&I3)|(I1&I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5613  */ #(
            .INIT(32'b10100010111100101111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5613  (
            .Z (_N10183_1044),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3&~I4)|(~I2&~I4)|(I2&~I3&I4)|(I0&I2&I3)|(I0&~I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5617  (
            .Z (_N10183_1048),
            .I0 (_N10183_1764),
            .I1 (_N10183_1765),
            .S (\u_lcd_rgb_char/bcd_data_y [3] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5618  (
            .Z (_N10183_1049),
            .I0 (_N10183_1766),
            .I1 (_N10183_1767),
            .S (\u_lcd_rgb_char/bcd_data_y [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5619  (
            .Z (_N10183_1050),
            .I0 (_N10183_1769),
            .I1 (_N10183_1768),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5621  */ #(
            .INIT(32'b11110011111011111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5621  (
            .Z (_N10183_1052),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I4)|(~I0&~I4)|(I0&~I1&I4)|(I1&~I3)|(~I0&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5625  */ #(
            .INIT(32'b10011011000100111001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5625  (
            .Z (_N10183_1056),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I2&~I4)|(~I1&~I2&I4)|(~I0&~I1&I4)|(~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_5626  */ #(
            .INIT(16'b1001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5626  (
            .Z (_N10183_1057),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5628  */ #(
            .INIT(32'b11111111110110111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5628  (
            .Z (_N10183_1059),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I4)|(I3&I4)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5629  */ #(
            .INIT(32'b11011111111011111110101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5629  (
            .Z (_N10183_1060),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(~I0&I3&I4)|(I1&~I3)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5630  */ #(
            .INIT(32'b11111011111011111110011111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5630  (
            .Z (_N10183_1061),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&I3&~I4)|(I1&~I3&I4)|(~I1&I3&I4)|(I0&I4)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5632  */ #(
            .INIT(32'b11111000000000000001111000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5632  (
            .Z (_N10183_1063),
            .I0 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&~I2&I3&~I4)|(I0&~I2&~I4)|(I2&I3&I4)|(I0&I1&~I2&I3)|(~I0&~I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5633  */ #(
            .INIT(32'b11111111110111111010101010001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5633  (
            .Z (_N10183_1064),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I4 (_N10183_1791));
	// LUT = (~I0&I4)|(I0&I3)|(I0&~I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5635  */ #(
            .INIT(32'b10101000101010000101001000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5635  (
            .Z (_N10183_1066),
            .I0 (_N10183_2782),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [2] ));
	// LUT = (ID&~I2&~I3&~I4)|(~ID&I2&I3&~I4)|(ID&~I1&~I2&~I4)|(I0&I2&I4)|(I0&I1&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5636  (
            .Z (_N10183_1067),
            .I0 (_N10183_1796),
            .I1 (_N10183_1795),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5638  */ #(
            .INIT(32'b10101011101110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5638  (
            .Z (_N10183_1069),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_1799));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(~I1&~I2&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5645  */ #(
            .INIT(32'b11100000000000000110001000010001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5645  (
            .Z (_N10183_1076),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I0&~I1&I3&~I4)|(I0&I2&I3&I4)|(~I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5646  */ #(
            .INIT(32'b10010001011101111110111100010111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5646  (
            .Z (_N10183_1077),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&I3&~I4)|(I0&I3&~I4)|(~I1&~I3&I4)|(~I0&~I3&I4)|(~I0&~I1&I4)|(~I1&~I2&~I3)|(~I0&~I2&~I3)|(~I0&~I1&~I3)|(I0&I1&I2&I3)|(~I0&~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5648  */ #(
            .INIT(32'b11111111001000000011111110100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5648  (
            .Z (_N10183_1079),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I0&I2&~I3&~I4)|(I3&I4)|(~I2&I3)|(~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5649  */ #(
            .INIT(32'b10111011000000010010000110111010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5649  (
            .Z (_N10183_1080),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&I2&~I3&~I4)|(I0&~I3&~I4)|(~I1&I3&I4)|(I0&I3&I4)|(~I0&~I1&~I2&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5653  (
            .Z (_N10183_1084),
            .I0 (_N10183_1822),
            .I1 (_N10183_1821),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5655  (
            .Z (_N10183_1086),
            .I0 (_N10183_1825),
            .I1 (_N10183_1826),
            .S (\u_lcd_rgb_char/bcd_data_x [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5656  (
            .Z (_N10183_1087),
            .I0 (_N10183_1827),
            .I1 (_N10183_1828),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5657  (
            .Z (_N10183_1088),
            .I0 (_N10183_1830),
            .I1 (_N10183_1829),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5658  (
            .Z (_N10183_1089),
            .I0 (_N10183_1832),
            .I1 (_N10183_1831),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5660  */ #(
            .INIT(32'b11111110111110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5660  (
            .Z (_N10183_1091),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1835));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5661  */ #(
            .INIT(32'b11101111111111111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5661  (
            .Z (_N10183_1092),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .ID (_N10183_1836));
	// LUT = (ID&~I4)|(~I3&I4)|(~I2&I4)|(I1&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5664  */ #(
            .INIT(32'b10111111110110011101101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5664  (
            .Z (_N10183_1095),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&I2&~I4)|(~I2&I3&I4)|(I0&I3&I4)|(~I0&I2&~I3)|(I0&~I2&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5665  */ #(
            .INIT(32'b10011000010110100111010011000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5665  (
            .Z (_N10183_1096),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&I2&~I3&~I4)|(~I1&I2&I3&~I4)|(~I0&I1&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(~I0&I1&I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5669  */ #(
            .INIT(32'b10111011111100111011101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5669  (
            .Z (_N10183_1100),
            .I0 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(I2&~I3)|(I0&I3)|(~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5671  */ #(
            .INIT(32'b10011111100111101111100111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5671  (
            .Z (_N10183_1102),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2&~I4)|(I1&~I2&I4)|(I0&~I2&I4)|(I1&~I2&~I3)|(I0&~I2&~I3)|(~I0&~I1&I3)|(~I0&~I1&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5674  */ #(
            .INIT(32'b11101000111111101110111111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5674  (
            .Z (_N10183_1105),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (_N10183_2852));
	// LUT = (~I2&~I4)|(ID&~I4)|(I2&~I3&I4)|(I0&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5677  */ #(
            .INIT(32'b11101100111011001101101110011011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5677  (
            .Z (_N10183_1108),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I2&~I4)|(~I0&~I1&~I4)|(I0&I2&I4)|(I1&I4)|(I1&I2&I3)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5683  */ #(
            .INIT(32'b11110111110001111101001111110011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5683  (
            .Z (_N10183_1114),
            .I0 (_N10183_2712),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .ID (_N10183_2642));
	// LUT = (~I1&~I3&~I4)|(~I1&I3&I4)|(~I0&I1&I4)|(~ID&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5685  */ #(
            .INIT(32'b11001100001100110000110100100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5685  (
            .Z (_N10183_1116),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I2&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I0&~I1&I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5686  */ #(
            .INIT(32'b11110110111111101111100010011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5686  (
            .Z (_N10183_1117),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I4)|(I0&~I1&I4)|(~I0&I1&I4)|(I0&I1&~I3)|(I2&I3)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5688  */ #(
            .INIT(32'b11101111011011110000100101101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5688  (
            .Z (_N10183_1119),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I0&I1&I4)|(I0&~I1&~I3)|(~I0&I1&~I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5690  */ #(
            .INIT(32'b10100101101001010001000100000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5690  (
            .Z (_N10183_1121),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I3&~I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5691_3  */ #(
            .INIT(32'b11001100000100011111111111111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5691_3  (
            .Z (_N10183_1122),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1004));
	// LUT = (I3&~I4)|(I2&~I4)|(I1&~I4)|(~ID&~I4)|(~I0&~I1&~I3&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5692  */ #(
            .INIT(32'b11110101000100010100010011110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5692  (
            .Z (_N10183_1123),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I2&~I3&~I4)|(~I0&I1&~I4)|(I2&I3&I4)|(~I0&~I1&I4)|(~I0&~I1&~I3)|(~I0&I1&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5695  (
            .Z (_N10183_1126),
            .I0 (_N10183_1884),
            .I1 (_N10183_1885),
            .S (\u_lcd_rgb_char/bcd_data_x [1] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5698  */ #(
            .INIT(32'b11111111101100110101100111101101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5698  (
            .Z (_N10183_1129),
            .I0 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(ID&~I1&I2&~I3)|(I0&ID&I2&~I3)|(ID&I1&~I2&I3)|(~ID&I2&I3)|(~ID&~I1&~I2)|(I0&~ID&I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5699  */ #(
            .INIT(32'b10101010101010101100111011001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5699  (
            .Z (_N10183_1130),
            .I0 (_N10183_1892),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [1] ));
	// LUT = (ID&~I2&I3&~I4)|(I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5701  */ #(
            .INIT(32'b11011110000100101101110000010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5701  (
            .Z (_N10183_1132),
            .I0 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I3 (_N10183_1894),
            .I4 (_N10183_1748),
            .ID (\u_lcd_rgb_char/bcd_data_x [0] ));
	// LUT = (~ID&~I1&I2&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5702  */ #(
            .INIT(32'b10101000011010000000001000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5702  (
            .Z (_N10183_1133),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&I1&I2&~I3&I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(I0&~I1&I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5704  */ #(
            .INIT(32'b10100101111100011110001001011010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5704  (
            .Z (_N10183_1135),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I3&~I4)|(I0&~I1&~I2&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&I2&I4)|(~I0&I2&~I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5705  */ #(
            .INIT(32'b11101010110010001100101010010100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5705  (
            .Z (_N10183_1136),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I0&I3&I4)|(I1&I2&I4)|(I0&I1&I4)|(I0&~I2&I3)|(I1&I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5706  */ #(
            .INIT(32'b10100010111100101111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5706  (
            .Z (_N10183_1137),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3&~I4)|(~I2&~I4)|(I2&~I3&I4)|(I0&I2&I3)|(I0&~I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5710  (
            .Z (_N10183_1141),
            .I0 (_N10183_1907),
            .I1 (_N10183_1908),
            .S (\u_lcd_rgb_char/bcd_data_x [3] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5711  (
            .Z (_N10183_1142),
            .I0 (_N10183_1909),
            .I1 (_N10183_1910),
            .S (\u_lcd_rgb_char/bcd_data_x [1] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5712  (
            .Z (_N10183_1143),
            .I0 (_N10183_1912),
            .I1 (_N10183_1911),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5714  */ #(
            .INIT(32'b11110011111011111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5714  (
            .Z (_N10183_1145),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I4)|(~I0&~I4)|(I0&~I1&I4)|(I1&~I3)|(~I0&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5717  */ #(
            .INIT(32'b10011011000100111001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5717  (
            .Z (_N10183_1148),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I2&~I4)|(~I1&~I2&I4)|(~I0&~I1&I4)|(~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_5718  */ #(
            .INIT(16'b1001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5718  (
            .Z (_N10183_1149),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5720  */ #(
            .INIT(32'b11111111110110111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5720  (
            .Z (_N10183_1151),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I4)|(I3&I4)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5721  */ #(
            .INIT(32'b11011111111011111110101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5721  (
            .Z (_N10183_1152),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(~I0&I3&I4)|(I1&~I3)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5722  */ #(
            .INIT(32'b11111011111011111110011111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5722  (
            .Z (_N10183_1153),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&I3&~I4)|(I1&~I3&I4)|(~I1&I3&I4)|(I0&I4)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5724  */ #(
            .INIT(32'b11111000000000000001111000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5724  (
            .Z (_N10183_1155),
            .I0 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&~I2&I3&~I4)|(I0&~I2&~I4)|(I2&I3&I4)|(I0&I1&~I2&I3)|(~I0&~I1&I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5726  */ #(
            .INIT(32'b10101000101010000101001000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5726  (
            .Z (_N10183_1157),
            .I0 (_N10183_2911),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [2] ));
	// LUT = (ID&~I2&~I3&~I4)|(~ID&I2&I3&~I4)|(ID&~I1&~I2&~I4)|(I0&I2&I4)|(I0&I1&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5727  (
            .Z (_N10183_1158),
            .I0 (_N10183_1936),
            .I1 (_N10183_1935),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5729  */ #(
            .INIT(32'b10101011101110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5729  (
            .Z (_N10183_1160),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_1938));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(~I1&~I2&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5736  */ #(
            .INIT(32'b11100000000000000110001000010001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5736  (
            .Z (_N10183_1167),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I0&~I1&I3&~I4)|(I0&I2&I3&I4)|(~I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5737  */ #(
            .INIT(32'b10010001011101111110111100010111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5737  (
            .Z (_N10183_1168),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&I3&~I4)|(I0&I3&~I4)|(~I1&~I3&I4)|(~I0&~I3&I4)|(~I0&~I1&I4)|(~I1&~I2&~I3)|(~I0&~I2&~I3)|(~I0&~I1&~I3)|(I0&I1&I2&I3)|(~I0&~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5739  */ #(
            .INIT(32'b11111111001000000011111110100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5739  (
            .Z (_N10183_1170),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I0&I2&~I3&~I4)|(I3&I4)|(~I2&I3)|(~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5740  */ #(
            .INIT(32'b10111011000000010010000110111010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5740  (
            .Z (_N10183_1171),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&I2&~I3&~I4)|(I0&~I3&~I4)|(~I1&I3&I4)|(I0&I3&I4)|(~I0&~I1&~I2&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5744  (
            .Z (_N10183_1175),
            .I0 (_N10183_1959),
            .I1 (_N10183_1958),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5746  (
            .Z (_N10183_1177),
            .I0 (_N10183_1962),
            .I1 (_N10183_1963),
            .S (\u_lcd_rgb_char/bcd_data_y [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5747  (
            .Z (_N10183_1178),
            .I0 (_N10183_1964),
            .I1 (_N10183_1965),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5748  (
            .Z (_N10183_1179),
            .I0 (_N10183_1967),
            .I1 (_N10183_1966),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5749  (
            .Z (_N10183_1180),
            .I0 (_N10183_1969),
            .I1 (_N10183_1968),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5751  */ #(
            .INIT(32'b11111110111110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5751  (
            .Z (_N10183_1182),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_1972));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5752  */ #(
            .INIT(32'b11101111111111111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5752  (
            .Z (_N10183_1183),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .ID (_N10183_1973));
	// LUT = (ID&~I4)|(~I3&I4)|(~I2&I4)|(I1&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5755  */ #(
            .INIT(32'b10111111110110011101101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5755  (
            .Z (_N10183_1186),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&I2&~I4)|(~I2&I3&I4)|(I0&I3&I4)|(~I0&I2&~I3)|(I0&~I2&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5756  */ #(
            .INIT(32'b10011000010110100111010011000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5756  (
            .Z (_N10183_1187),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&I2&~I3&~I4)|(~I1&I2&I3&~I4)|(~I0&I1&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(~I0&I1&I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5760  */ #(
            .INIT(32'b10111011111100111011101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5760  (
            .Z (_N10183_1191),
            .I0 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(I2&~I3)|(I0&I3)|(~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5762  */ #(
            .INIT(32'b10011111100111101111100111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5762  (
            .Z (_N10183_1193),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2&~I4)|(I1&~I2&I4)|(I0&~I2&I4)|(I1&~I2&~I3)|(I0&~I2&~I3)|(~I0&~I1&I3)|(~I0&~I1&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5765  */ #(
            .INIT(32'b11101000111111101110111111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5765  (
            .Z (_N10183_1196),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (_N10183_2976));
	// LUT = (~I2&~I4)|(ID&~I4)|(I2&~I3&I4)|(I0&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5768  */ #(
            .INIT(32'b11101100111011001101101110011011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5768  (
            .Z (_N10183_1199),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I2&~I4)|(~I0&~I1&~I4)|(I0&I2&I4)|(I1&I4)|(I1&I2&I3)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5774  */ #(
            .INIT(32'b11110111110001111101001111110011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5774  (
            .Z (_N10183_1205),
            .I0 (_N10183_2712),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .ID (_N10183_2642));
	// LUT = (~I1&~I3&~I4)|(~I1&I3&I4)|(~I0&I1&I4)|(~ID&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5776  */ #(
            .INIT(32'b11001100001100110000110100100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5776  (
            .Z (_N10183_1207),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I2&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I0&~I1&I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5777  */ #(
            .INIT(32'b11110110111111101111100010011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5777  (
            .Z (_N10183_1208),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I4)|(I0&~I1&I4)|(~I0&I1&I4)|(I0&I1&~I3)|(I2&I3)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5779  */ #(
            .INIT(32'b11101111011011110000100101101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5779  (
            .Z (_N10183_1210),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I0&I1&I4)|(I0&~I1&~I3)|(~I0&I1&~I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5781  */ #(
            .INIT(32'b10100101101001010001000100000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5781  (
            .Z (_N10183_1212),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I3&~I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5782_3  */ #(
            .INIT(32'b11001100000100011111111111111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5782_3  (
            .Z (_N10183_1213),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1004));
	// LUT = (I3&~I4)|(I2&~I4)|(I1&~I4)|(~ID&~I4)|(~I0&~I1&~I3&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5783  */ #(
            .INIT(32'b11110101000100010100010011110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5783  (
            .Z (_N10183_1214),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I2&~I3&~I4)|(~I0&I1&~I4)|(I2&I3&I4)|(~I0&~I1&I4)|(~I0&~I1&~I3)|(~I0&I1&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5786  (
            .Z (_N10183_1217),
            .I0 (_N10183_2021),
            .I1 (_N10183_2022),
            .S (\u_lcd_rgb_char/bcd_data_y [5] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5789  */ #(
            .INIT(32'b11111111101100110101100111101101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5789  (
            .Z (_N10183_1220),
            .I0 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(ID&~I1&I2&~I3)|(I0&ID&I2&~I3)|(ID&I1&~I2&I3)|(~ID&I2&I3)|(~ID&~I1&~I2)|(I0&~ID&I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5790  */ #(
            .INIT(32'b10101010101010101100111011001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5790  (
            .Z (_N10183_1221),
            .I0 (_N10183_2029),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [5] ));
	// LUT = (ID&~I2&I3&~I4)|(I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5792  */ #(
            .INIT(32'b11011110000100101101110000010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5792  (
            .Z (_N10183_1223),
            .I0 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I3 (_N10183_2031),
            .I4 (_N10183_1748),
            .ID (\u_lcd_rgb_char/bcd_data_y [4] ));
	// LUT = (~ID&~I1&I2&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5793  */ #(
            .INIT(32'b10101000011010000000001000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5793  (
            .Z (_N10183_1224),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&I1&I2&~I3&I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(I0&~I1&I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5795  */ #(
            .INIT(32'b10100101111100011110001001011010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5795  (
            .Z (_N10183_1226),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I3&~I4)|(I0&~I1&~I2&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&I2&I4)|(~I0&I2&~I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5796  */ #(
            .INIT(32'b11101010110010001100101010010100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5796  (
            .Z (_N10183_1227),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I0&I3&I4)|(I1&I2&I4)|(I0&I1&I4)|(I0&~I2&I3)|(I1&I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5797  */ #(
            .INIT(32'b10100010111100101111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5797  (
            .Z (_N10183_1228),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3&~I4)|(~I2&~I4)|(I2&~I3&I4)|(I0&I2&I3)|(I0&~I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5801  (
            .Z (_N10183_1232),
            .I0 (_N10183_2044),
            .I1 (_N10183_2045),
            .S (\u_lcd_rgb_char/bcd_data_y [7] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5802  (
            .Z (_N10183_1233),
            .I0 (_N10183_2046),
            .I1 (_N10183_2047),
            .S (\u_lcd_rgb_char/bcd_data_y [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5803  (
            .Z (_N10183_1234),
            .I0 (_N10183_2049),
            .I1 (_N10183_2048),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5805  */ #(
            .INIT(32'b11110011111011111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5805  (
            .Z (_N10183_1236),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I4)|(~I0&~I4)|(I0&~I1&I4)|(I1&~I3)|(~I0&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5808  */ #(
            .INIT(32'b10011011000100111001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5808  (
            .Z (_N10183_1239),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I2&~I4)|(~I1&~I2&I4)|(~I0&~I1&I4)|(~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_5809  */ #(
            .INIT(16'b1001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5809  (
            .Z (_N10183_1240),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5811  */ #(
            .INIT(32'b11111111110110111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5811  (
            .Z (_N10183_1242),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I4)|(I3&I4)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5812  */ #(
            .INIT(32'b11011111111011111110101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5812  (
            .Z (_N10183_1243),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(~I0&I3&I4)|(I1&~I3)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5813  */ #(
            .INIT(32'b11111011111011111110011111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5813  (
            .Z (_N10183_1244),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&I3&~I4)|(I1&~I3&I4)|(~I1&I3&I4)|(I0&I4)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5815  */ #(
            .INIT(32'b11111000000000000001111000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5815  (
            .Z (_N10183_1246),
            .I0 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&~I2&I3&~I4)|(I0&~I2&~I4)|(I2&I3&I4)|(I0&I1&~I2&I3)|(~I0&~I1&I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5817  */ #(
            .INIT(32'b10101000101010000101001000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5817  (
            .Z (_N10183_1248),
            .I0 (_N10183_3032),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [6] ));
	// LUT = (ID&~I2&~I3&~I4)|(~ID&I2&I3&~I4)|(ID&~I1&~I2&~I4)|(I0&I2&I4)|(I0&I1&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5818  (
            .Z (_N10183_1249),
            .I0 (_N10183_2073),
            .I1 (_N10183_2072),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5820  */ #(
            .INIT(32'b10101011101110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5820  (
            .Z (_N10183_1251),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_2075));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(~I1&~I2&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5827  */ #(
            .INIT(32'b11100000000000000110001000010001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5827  (
            .Z (_N10183_1258),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I0&~I1&I3&~I4)|(I0&I2&I3&I4)|(~I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5828  */ #(
            .INIT(32'b10010001011101111110111100010111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5828  (
            .Z (_N10183_1259),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&I3&~I4)|(I0&I3&~I4)|(~I1&~I3&I4)|(~I0&~I3&I4)|(~I0&~I1&I4)|(~I1&~I2&~I3)|(~I0&~I2&~I3)|(~I0&~I1&~I3)|(I0&I1&I2&I3)|(~I0&~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5830  */ #(
            .INIT(32'b11111111001000000011111110100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5830  (
            .Z (_N10183_1261),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I0&I2&~I3&~I4)|(I3&I4)|(~I2&I3)|(~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5831  */ #(
            .INIT(32'b10111011000000010010000110111010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5831  (
            .Z (_N10183_1262),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&I2&~I3&~I4)|(I0&~I3&~I4)|(~I1&I3&I4)|(I0&I3&I4)|(~I0&~I1&~I2&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5835  (
            .Z (_N10183_1266),
            .I0 (_N10183_2096),
            .I1 (_N10183_2095),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5837  (
            .Z (_N10183_1268),
            .I0 (_N10183_2099),
            .I1 (_N10183_2100),
            .S (\u_lcd_rgb_char/bcd_data_x [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5838  (
            .Z (_N10183_1269),
            .I0 (_N10183_2101),
            .I1 (_N10183_2102),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5839  (
            .Z (_N10183_1270),
            .I0 (_N10183_2104),
            .I1 (_N10183_2103),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5840  (
            .Z (_N10183_1271),
            .I0 (_N10183_2106),
            .I1 (_N10183_2105),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5842  */ #(
            .INIT(32'b11111110111110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5842  (
            .Z (_N10183_1273),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_2109));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5843  */ #(
            .INIT(32'b11101111111111111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5843  (
            .Z (_N10183_1274),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .ID (_N10183_2110));
	// LUT = (ID&~I4)|(~I3&I4)|(~I2&I4)|(I1&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5846  */ #(
            .INIT(32'b10111111110110011101101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5846  (
            .Z (_N10183_1277),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&I2&~I4)|(~I2&I3&I4)|(I0&I3&I4)|(~I0&I2&~I3)|(I0&~I2&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5847  */ #(
            .INIT(32'b10011000010110100111010011000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5847  (
            .Z (_N10183_1278),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&I2&~I3&~I4)|(~I1&I2&I3&~I4)|(~I0&I1&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(~I0&I1&I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5851  */ #(
            .INIT(32'b10111011111100111011101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5851  (
            .Z (_N10183_1282),
            .I0 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(I2&~I3)|(I0&I3)|(~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5853  */ #(
            .INIT(32'b10011111100111101111100111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5853  (
            .Z (_N10183_1284),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2&~I4)|(I1&~I2&I4)|(I0&~I2&I4)|(I1&~I2&~I3)|(I0&~I2&~I3)|(~I0&~I1&I3)|(~I0&~I1&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5856  */ #(
            .INIT(32'b11101000111111101110111111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5856  (
            .Z (_N10183_1287),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (_N10183_3097));
	// LUT = (~I2&~I4)|(ID&~I4)|(I2&~I3&I4)|(I0&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5859  */ #(
            .INIT(32'b11101100111011001101101110011011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5859  (
            .Z (_N10183_1290),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I2&~I4)|(~I0&~I1&~I4)|(I0&I2&I4)|(I1&I4)|(I1&I2&I3)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5865  */ #(
            .INIT(32'b11110111110001111101001111110011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5865  (
            .Z (_N10183_1296),
            .I0 (_N10183_2712),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .ID (_N10183_2642));
	// LUT = (~I1&~I3&~I4)|(~I1&I3&I4)|(~I0&I1&I4)|(~ID&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5867  */ #(
            .INIT(32'b11001100001100110000110100100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5867  (
            .Z (_N10183_1298),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I2&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I0&~I1&I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5868  */ #(
            .INIT(32'b11110110111111101111100010011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5868  (
            .Z (_N10183_1299),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I4)|(I0&~I1&I4)|(~I0&I1&I4)|(I0&I1&~I3)|(I2&I3)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5870  */ #(
            .INIT(32'b11101111011011110000100101101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5870  (
            .Z (_N10183_1301),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I0&I1&I4)|(I0&~I1&~I3)|(~I0&I1&~I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5872  */ #(
            .INIT(32'b10100101101001010001000100000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5872  (
            .Z (_N10183_1303),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I3&~I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5873_3  */ #(
            .INIT(32'b11001100000100011111111111111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5873_3  (
            .Z (_N10183_1304),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1004));
	// LUT = (I3&~I4)|(I2&~I4)|(I1&~I4)|(~ID&~I4)|(~I0&~I1&~I3&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5874  */ #(
            .INIT(32'b11110101000100010100010011110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5874  (
            .Z (_N10183_1305),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I2&~I3&~I4)|(~I0&I1&~I4)|(I2&I3&I4)|(~I0&~I1&I4)|(~I0&~I1&~I3)|(~I0&I1&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5877  (
            .Z (_N10183_1308),
            .I0 (_N10183_2158),
            .I1 (_N10183_2159),
            .S (\u_lcd_rgb_char/bcd_data_x [5] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5880  */ #(
            .INIT(32'b11111111101100110101100111101101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5880  (
            .Z (_N10183_1311),
            .I0 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(ID&~I1&I2&~I3)|(I0&ID&I2&~I3)|(ID&I1&~I2&I3)|(~ID&I2&I3)|(~ID&~I1&~I2)|(I0&~ID&I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5881  */ #(
            .INIT(32'b10101010101010101100111011001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5881  (
            .Z (_N10183_1312),
            .I0 (_N10183_2166),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [5] ));
	// LUT = (ID&~I2&I3&~I4)|(I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5883  */ #(
            .INIT(32'b11011110000100101101110000010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5883  (
            .Z (_N10183_1314),
            .I0 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I3 (_N10183_2168),
            .I4 (_N10183_1748),
            .ID (\u_lcd_rgb_char/bcd_data_x [4] ));
	// LUT = (~ID&~I1&I2&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5884  */ #(
            .INIT(32'b10101000011010000000001000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5884  (
            .Z (_N10183_1315),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&I1&I2&~I3&I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(I0&~I1&I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5886  */ #(
            .INIT(32'b10100101111100011110001001011010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5886  (
            .Z (_N10183_1317),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I3&~I4)|(I0&~I1&~I2&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&I2&I4)|(~I0&I2&~I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5887  */ #(
            .INIT(32'b11101010110010001100101010010100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5887  (
            .Z (_N10183_1318),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I0&I3&I4)|(I1&I2&I4)|(I0&I1&I4)|(I0&~I2&I3)|(I1&I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5888  */ #(
            .INIT(32'b10100010111100101111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5888  (
            .Z (_N10183_1319),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3&~I4)|(~I2&~I4)|(I2&~I3&I4)|(I0&I2&I3)|(I0&~I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5892  (
            .Z (_N10183_1323),
            .I0 (_N10183_2181),
            .I1 (_N10183_2182),
            .S (\u_lcd_rgb_char/bcd_data_x [7] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5893  (
            .Z (_N10183_1324),
            .I0 (_N10183_2183),
            .I1 (_N10183_2184),
            .S (\u_lcd_rgb_char/bcd_data_x [5] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5894  (
            .Z (_N10183_1325),
            .I0 (_N10183_2186),
            .I1 (_N10183_2185),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5896  */ #(
            .INIT(32'b11110011111011111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5896  (
            .Z (_N10183_1327),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I4)|(~I0&~I4)|(I0&~I1&I4)|(I1&~I3)|(~I0&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5899  */ #(
            .INIT(32'b10011011000100111001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5899  (
            .Z (_N10183_1330),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I2&~I4)|(~I1&~I2&I4)|(~I0&~I1&I4)|(~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_5900  */ #(
            .INIT(16'b1001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5900  (
            .Z (_N10183_1331),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5902  */ #(
            .INIT(32'b11111111110110111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5902  (
            .Z (_N10183_1333),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I4)|(I3&I4)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5903  */ #(
            .INIT(32'b11011111111011111110101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5903  (
            .Z (_N10183_1334),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(~I0&I3&I4)|(I1&~I3)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5904  */ #(
            .INIT(32'b11111011111011111110011111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5904  (
            .Z (_N10183_1335),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&I3&~I4)|(I1&~I3&I4)|(~I1&I3&I4)|(I0&I4)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5906  */ #(
            .INIT(32'b11111000000000000001111000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5906  (
            .Z (_N10183_1337),
            .I0 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&~I2&I3&~I4)|(I0&~I2&~I4)|(I2&I3&I4)|(I0&I1&~I2&I3)|(~I0&~I1&I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5908  */ #(
            .INIT(32'b10101000101010000101001000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5908  (
            .Z (_N10183_1339),
            .I0 (_N10183_3153),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [6] ));
	// LUT = (ID&~I2&~I3&~I4)|(~ID&I2&I3&~I4)|(ID&~I1&~I2&~I4)|(I0&I2&I4)|(I0&I1&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5909  (
            .Z (_N10183_1340),
            .I0 (_N10183_2210),
            .I1 (_N10183_2209),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5911  */ #(
            .INIT(32'b10101011101110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5911  (
            .Z (_N10183_1342),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_2212));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(~I1&~I2&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5918  */ #(
            .INIT(32'b11100000000000000110001000010001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5918  (
            .Z (_N10183_1349),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I0&~I1&I3&~I4)|(I0&I2&I3&I4)|(~I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5919  */ #(
            .INIT(32'b10010001011101111110111100010111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5919  (
            .Z (_N10183_1350),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&I3&~I4)|(I0&I3&~I4)|(~I1&~I3&I4)|(~I0&~I3&I4)|(~I0&~I1&I4)|(~I1&~I2&~I3)|(~I0&~I2&~I3)|(~I0&~I1&~I3)|(I0&I1&I2&I3)|(~I0&~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5921  */ #(
            .INIT(32'b11111111001000000011111110100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5921  (
            .Z (_N10183_1352),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I0&I2&~I3&~I4)|(I3&I4)|(~I2&I3)|(~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5922  */ #(
            .INIT(32'b10111011000000010010000110111010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5922  (
            .Z (_N10183_1353),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&I2&~I3&~I4)|(I0&~I3&~I4)|(~I1&I3&I4)|(I0&I3&I4)|(~I0&~I1&~I2&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5926  (
            .Z (_N10183_1357),
            .I0 (_N10183_2233),
            .I1 (_N10183_2232),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5928  (
            .Z (_N10183_1359),
            .I0 (_N10183_2236),
            .I1 (_N10183_2237),
            .S (\u_lcd_rgb_char/bcd_data_y [9] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5929  (
            .Z (_N10183_1360),
            .I0 (_N10183_2238),
            .I1 (_N10183_2239),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5930  (
            .Z (_N10183_1361),
            .I0 (_N10183_2241),
            .I1 (_N10183_2240),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5931  (
            .Z (_N10183_1362),
            .I0 (_N10183_2243),
            .I1 (_N10183_2242),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5933  */ #(
            .INIT(32'b11111110111110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5933  (
            .Z (_N10183_1364),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_2246));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5934  */ #(
            .INIT(32'b11101111111111111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5934  (
            .Z (_N10183_1365),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .ID (_N10183_2247));
	// LUT = (ID&~I4)|(~I3&I4)|(~I2&I4)|(I1&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5937  */ #(
            .INIT(32'b10111111110110011101101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5937  (
            .Z (_N10183_1368),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&I2&~I4)|(~I2&I3&I4)|(I0&I3&I4)|(~I0&I2&~I3)|(I0&~I2&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5938  */ #(
            .INIT(32'b10011000010110100111010011000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5938  (
            .Z (_N10183_1369),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&I2&~I3&~I4)|(~I1&I2&I3&~I4)|(~I0&I1&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(~I0&I1&I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5942  */ #(
            .INIT(32'b10111011111100111011101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5942  (
            .Z (_N10183_1373),
            .I0 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(I2&~I3)|(I0&I3)|(~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5944  */ #(
            .INIT(32'b10011111100111101111100111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_5944  (
            .Z (_N10183_1375),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2&~I4)|(I1&~I2&I4)|(I0&~I2&I4)|(I1&~I2&~I3)|(I0&~I2&~I3)|(~I0&~I1&I3)|(~I0&~I1&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5947  */ #(
            .INIT(32'b11101000111111101110111111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5947  (
            .Z (_N10183_1378),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (_N10183_3218));
	// LUT = (~I2&~I4)|(ID&~I4)|(I2&~I3&I4)|(I0&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5950  */ #(
            .INIT(32'b11101100111011001101101110011011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5950  (
            .Z (_N10183_1381),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I2&~I4)|(~I0&~I1&~I4)|(I0&I2&I4)|(I1&I4)|(I1&I2&I3)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5956  */ #(
            .INIT(32'b11110111110001111101001111110011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5956  (
            .Z (_N10183_1387),
            .I0 (_N10183_2712),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .ID (_N10183_2642));
	// LUT = (~I1&~I3&~I4)|(~I1&I3&I4)|(~I0&I1&I4)|(~ID&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5958  */ #(
            .INIT(32'b11001100001100110000110100100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5958  (
            .Z (_N10183_1389),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I2&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I0&~I1&I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5959  */ #(
            .INIT(32'b11110110111111101111100010011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5959  (
            .Z (_N10183_1390),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I4)|(I0&~I1&I4)|(~I0&I1&I4)|(I0&I1&~I3)|(I2&I3)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5961  */ #(
            .INIT(32'b11101111011011110000100101101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5961  (
            .Z (_N10183_1392),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I0&I1&I4)|(I0&~I1&~I3)|(~I0&I1&~I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5963  */ #(
            .INIT(32'b10100101101001010001000100000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5963  (
            .Z (_N10183_1394),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I3&~I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5964_3  */ #(
            .INIT(32'b11001100000100011111111111111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5964_3  (
            .Z (_N10183_1395),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1004));
	// LUT = (I3&~I4)|(I2&~I4)|(I1&~I4)|(~ID&~I4)|(~I0&~I1&~I3&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5965  */ #(
            .INIT(32'b11110101000100010100010011110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5965  (
            .Z (_N10183_1396),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I2&~I3&~I4)|(~I0&I1&~I4)|(I2&I3&I4)|(~I0&~I1&I4)|(~I0&~I1&~I3)|(~I0&I1&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5968  (
            .Z (_N10183_1399),
            .I0 (_N10183_2295),
            .I1 (_N10183_2296),
            .S (\u_lcd_rgb_char/bcd_data_y [9] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5971  */ #(
            .INIT(32'b11111111101100110101100111101101))
        \u_lcd_rgb_char/u_lcd_display/N9971_5971  (
            .Z (_N10183_1402),
            .I0 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(ID&~I1&I2&~I3)|(I0&ID&I2&~I3)|(ID&I1&~I2&I3)|(~ID&I2&I3)|(~ID&~I1&~I2)|(I0&~ID&I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5972  */ #(
            .INIT(32'b10101010101010101100111011001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5972  (
            .Z (_N10183_1403),
            .I0 (_N10183_2303),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [9] ));
	// LUT = (ID&~I2&I3&~I4)|(I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5974  */ #(
            .INIT(32'b11011110000100101101110000010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5974  (
            .Z (_N10183_1405),
            .I0 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I3 (_N10183_2305),
            .I4 (_N10183_1748),
            .ID (\u_lcd_rgb_char/bcd_data_y [8] ));
	// LUT = (~ID&~I1&I2&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5975  */ #(
            .INIT(32'b10101000011010000000001000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_5975  (
            .Z (_N10183_1406),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&I1&I2&~I3&I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(I0&~I1&I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5977  */ #(
            .INIT(32'b10100101111100011110001001011010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5977  (
            .Z (_N10183_1408),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I3&~I4)|(I0&~I1&~I2&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&I2&I4)|(~I0&I2&~I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5978  */ #(
            .INIT(32'b11101010110010001100101010010100))
        \u_lcd_rgb_char/u_lcd_display/N9971_5978  (
            .Z (_N10183_1409),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I0&I3&I4)|(I1&I2&I4)|(I0&I1&I4)|(I0&~I2&I3)|(I1&I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5979  */ #(
            .INIT(32'b10100010111100101111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5979  (
            .Z (_N10183_1410),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3&~I4)|(~I2&~I4)|(I2&~I3&I4)|(I0&I2&I3)|(I0&~I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5983  (
            .Z (_N10183_1414),
            .I0 (_N10183_2318),
            .I1 (_N10183_2319),
            .S (\u_lcd_rgb_char/bcd_data_y [11] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5984  (
            .Z (_N10183_1415),
            .I0 (_N10183_2320),
            .I1 (_N10183_2321),
            .S (\u_lcd_rgb_char/bcd_data_y [9] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_5985  (
            .Z (_N10183_1416),
            .I0 (_N10183_2323),
            .I1 (_N10183_2322),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5987  */ #(
            .INIT(32'b11110011111011111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5987  (
            .Z (_N10183_1418),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I4)|(~I0&~I4)|(I0&~I1&I4)|(I1&~I3)|(~I0&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5990  */ #(
            .INIT(32'b10011011000100111001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5990  (
            .Z (_N10183_1421),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I2&~I4)|(~I1&~I2&I4)|(~I0&~I1&I4)|(~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_5991  */ #(
            .INIT(16'b1001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_5991  (
            .Z (_N10183_1422),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5993  */ #(
            .INIT(32'b11111111110110111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5993  (
            .Z (_N10183_1424),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I4)|(I3&I4)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5994  */ #(
            .INIT(32'b11011111111011111110101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_5994  (
            .Z (_N10183_1425),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(~I0&I3&I4)|(I1&~I3)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5995  */ #(
            .INIT(32'b11111011111011111110011111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_5995  (
            .Z (_N10183_1426),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&I3&~I4)|(I1&~I3&I4)|(~I1&I3&I4)|(I0&I4)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_5997  */ #(
            .INIT(32'b11111000000000000001111000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5997  (
            .Z (_N10183_1428),
            .I0 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&~I2&I3&~I4)|(I0&~I2&~I4)|(I2&I3&I4)|(I0&I1&~I2&I3)|(~I0&~I1&I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_5999  */ #(
            .INIT(32'b10101000101010000101001000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_5999  (
            .Z (_N10183_1430),
            .I0 (_N10183_3274),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_y [10] ));
	// LUT = (ID&~I2&~I3&~I4)|(~ID&I2&I3&~I4)|(ID&~I1&~I2&~I4)|(I0&I2&I4)|(I0&I1&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6000  (
            .Z (_N10183_1431),
            .I0 (_N10183_2347),
            .I1 (_N10183_2346),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6002  */ #(
            .INIT(32'b10101011101110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6002  (
            .Z (_N10183_1433),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_2349));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(~I1&~I2&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6009  */ #(
            .INIT(32'b11100000000000000110001000010001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6009  (
            .Z (_N10183_1440),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I0&~I1&I3&~I4)|(I0&I2&I3&I4)|(~I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6010  */ #(
            .INIT(32'b10010001011101111110111100010111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6010  (
            .Z (_N10183_1441),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&I3&~I4)|(I0&I3&~I4)|(~I1&~I3&I4)|(~I0&~I3&I4)|(~I0&~I1&I4)|(~I1&~I2&~I3)|(~I0&~I2&~I3)|(~I0&~I1&~I3)|(I0&I1&I2&I3)|(~I0&~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6012  */ #(
            .INIT(32'b11111111001000000011111110100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6012  (
            .Z (_N10183_1443),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I0&I2&~I3&~I4)|(I3&I4)|(~I2&I3)|(~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6013  */ #(
            .INIT(32'b10111011000000010010000110111010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6013  (
            .Z (_N10183_1444),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&I2&~I3&~I4)|(I0&~I3&~I4)|(~I1&I3&I4)|(I0&I3&I4)|(~I0&~I1&~I2&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6017  (
            .Z (_N10183_1448),
            .I0 (_N10183_2370),
            .I1 (_N10183_2369),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6019  (
            .Z (_N10183_1450),
            .I0 (_N10183_2373),
            .I1 (_N10183_2374),
            .S (\u_lcd_rgb_char/bcd_data_x [9] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6020  (
            .Z (_N10183_1451),
            .I0 (_N10183_2375),
            .I1 (_N10183_2376),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6021  (
            .Z (_N10183_1452),
            .I0 (_N10183_2378),
            .I1 (_N10183_2377),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6022  (
            .Z (_N10183_1453),
            .I0 (_N10183_2380),
            .I1 (_N10183_2379),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6024  */ #(
            .INIT(32'b11111110111110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6024  (
            .Z (_N10183_1455),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_2383));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6025  */ #(
            .INIT(32'b11101111111111111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6025  (
            .Z (_N10183_1456),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .ID (_N10183_2384));
	// LUT = (ID&~I4)|(~I3&I4)|(~I2&I4)|(I1&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6028  */ #(
            .INIT(32'b10111111110110011101101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6028  (
            .Z (_N10183_1459),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&I2&~I4)|(~I2&I3&I4)|(I0&I3&I4)|(~I0&I2&~I3)|(I0&~I2&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6029  */ #(
            .INIT(32'b10011000010110100111010011000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6029  (
            .Z (_N10183_1460),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&I2&~I3&~I4)|(~I1&I2&I3&~I4)|(~I0&I1&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(~I0&I1&I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6033  */ #(
            .INIT(32'b10111011111100111011101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6033  (
            .Z (_N10183_1464),
            .I0 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(I2&~I3)|(I0&I3)|(~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6035  */ #(
            .INIT(32'b10011111100111101111100111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6035  (
            .Z (_N10183_1466),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2&~I4)|(I1&~I2&I4)|(I0&~I2&I4)|(I1&~I2&~I3)|(I0&~I2&~I3)|(~I0&~I1&I3)|(~I0&~I1&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6038  */ #(
            .INIT(32'b11101000111111101110111111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6038  (
            .Z (_N10183_1469),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (_N10183_3339));
	// LUT = (~I2&~I4)|(ID&~I4)|(I2&~I3&I4)|(I0&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6041  */ #(
            .INIT(32'b11101100111011001101101110011011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6041  (
            .Z (_N10183_1472),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I2&~I4)|(~I0&~I1&~I4)|(I0&I2&I4)|(I1&I4)|(I1&I2&I3)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6047  */ #(
            .INIT(32'b11110111110001111101001111110011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6047  (
            .Z (_N10183_1478),
            .I0 (_N10183_2712),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .ID (_N10183_2642));
	// LUT = (~I1&~I3&~I4)|(~I1&I3&I4)|(~I0&I1&I4)|(~ID&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6049  */ #(
            .INIT(32'b11001100001100110000110100100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6049  (
            .Z (_N10183_1480),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I2&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I0&~I1&I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6050  */ #(
            .INIT(32'b11110110111111101111100010011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6050  (
            .Z (_N10183_1481),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I4)|(I0&~I1&I4)|(~I0&I1&I4)|(I0&I1&~I3)|(I2&I3)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6052  */ #(
            .INIT(32'b11101111011011110000100101101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6052  (
            .Z (_N10183_1483),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I0&I1&I4)|(I0&~I1&~I3)|(~I0&I1&~I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6054  */ #(
            .INIT(32'b10100101101001010001000100000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6054  (
            .Z (_N10183_1485),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I3&~I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6055_3  */ #(
            .INIT(32'b11001100000100011111111111111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6055_3  (
            .Z (_N10183_1486),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1004));
	// LUT = (I3&~I4)|(I2&~I4)|(I1&~I4)|(~ID&~I4)|(~I0&~I1&~I3&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6056  */ #(
            .INIT(32'b11110101000100010100010011110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6056  (
            .Z (_N10183_1487),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I2&~I3&~I4)|(~I0&I1&~I4)|(I2&I3&I4)|(~I0&~I1&I4)|(~I0&~I1&~I3)|(~I0&I1&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6059  (
            .Z (_N10183_1490),
            .I0 (_N10183_2432),
            .I1 (_N10183_2433),
            .S (\u_lcd_rgb_char/bcd_data_x [9] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6062  */ #(
            .INIT(32'b11111111101100110101100111101101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6062  (
            .Z (_N10183_1493),
            .I0 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(ID&~I1&I2&~I3)|(I0&ID&I2&~I3)|(ID&I1&~I2&I3)|(~ID&I2&I3)|(~ID&~I1&~I2)|(I0&~ID&I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6063  */ #(
            .INIT(32'b10101010101010101100111011001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6063  (
            .Z (_N10183_1494),
            .I0 (_N10183_2440),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [9] ));
	// LUT = (ID&~I2&I3&~I4)|(I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6065  */ #(
            .INIT(32'b11011110000100101101110000010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6065  (
            .Z (_N10183_1496),
            .I0 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I3 (_N10183_2442),
            .I4 (_N10183_1748),
            .ID (\u_lcd_rgb_char/bcd_data_x [8] ));
	// LUT = (~ID&~I1&I2&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6066  */ #(
            .INIT(32'b10101000011010000000001000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6066  (
            .Z (_N10183_1497),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&I1&I2&~I3&I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(I0&~I1&I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6068  */ #(
            .INIT(32'b10100101111100011110001001011010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6068  (
            .Z (_N10183_1499),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I3&~I4)|(I0&~I1&~I2&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&I2&I4)|(~I0&I2&~I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6069  */ #(
            .INIT(32'b11101010110010001100101010010100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6069  (
            .Z (_N10183_1500),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I0&I3&I4)|(I1&I2&I4)|(I0&I1&I4)|(I0&~I2&I3)|(I1&I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6070  */ #(
            .INIT(32'b10100010111100101111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6070  (
            .Z (_N10183_1501),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3&~I4)|(~I2&~I4)|(I2&~I3&I4)|(I0&I2&I3)|(I0&~I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6074  (
            .Z (_N10183_1505),
            .I0 (_N10183_2455),
            .I1 (_N10183_2456),
            .S (\u_lcd_rgb_char/bcd_data_x [11] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6075  (
            .Z (_N10183_1506),
            .I0 (_N10183_2457),
            .I1 (_N10183_2458),
            .S (\u_lcd_rgb_char/bcd_data_x [9] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6076  (
            .Z (_N10183_1507),
            .I0 (_N10183_2460),
            .I1 (_N10183_2459),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6078  */ #(
            .INIT(32'b11110011111011111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6078  (
            .Z (_N10183_1509),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I4)|(~I0&~I4)|(I0&~I1&I4)|(I1&~I3)|(~I0&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6081  */ #(
            .INIT(32'b10011011000100111001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6081  (
            .Z (_N10183_1512),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I2&~I4)|(~I1&~I2&I4)|(~I0&~I1&I4)|(~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6082  */ #(
            .INIT(16'b1001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6082  (
            .Z (_N10183_1513),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6084  */ #(
            .INIT(32'b11111111110110111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6084  (
            .Z (_N10183_1515),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I4)|(I3&I4)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6085  */ #(
            .INIT(32'b11011111111011111110101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6085  (
            .Z (_N10183_1516),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(~I0&I3&I4)|(I1&~I3)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6086  */ #(
            .INIT(32'b11111011111011111110011111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6086  (
            .Z (_N10183_1517),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&I3&~I4)|(I1&~I3&I4)|(~I1&I3&I4)|(I0&I4)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6088  */ #(
            .INIT(32'b11111000000000000001111000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6088  (
            .Z (_N10183_1519),
            .I0 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&~I2&I3&~I4)|(I0&~I2&~I4)|(I2&I3&I4)|(I0&I1&~I2&I3)|(~I0&~I1&I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6090  */ #(
            .INIT(32'b10101000101010000101001000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6090  (
            .Z (_N10183_1521),
            .I0 (_N10183_3395),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [10] ));
	// LUT = (ID&~I2&~I3&~I4)|(~ID&I2&I3&~I4)|(ID&~I1&~I2&~I4)|(I0&I2&I4)|(I0&I1&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6091  (
            .Z (_N10183_1522),
            .I0 (_N10183_2484),
            .I1 (_N10183_2483),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6093  */ #(
            .INIT(32'b10101011101110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6093  (
            .Z (_N10183_1524),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_2486));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(~I1&~I2&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6100  */ #(
            .INIT(32'b11100000000000000110001000010001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6100  (
            .Z (_N10183_1531),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I0&~I1&I3&~I4)|(I0&I2&I3&I4)|(~I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6101  */ #(
            .INIT(32'b10010001011101111110111100010111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6101  (
            .Z (_N10183_1532),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&I3&~I4)|(I0&I3&~I4)|(~I1&~I3&I4)|(~I0&~I3&I4)|(~I0&~I1&I4)|(~I1&~I2&~I3)|(~I0&~I2&~I3)|(~I0&~I1&~I3)|(I0&I1&I2&I3)|(~I0&~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6103  */ #(
            .INIT(32'b11111111001000000011111110100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6103  (
            .Z (_N10183_1534),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I0&I2&~I3&~I4)|(I3&I4)|(~I2&I3)|(~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6104  */ #(
            .INIT(32'b10111011000000010010000110111010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6104  (
            .Z (_N10183_1535),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&I2&~I3&~I4)|(I0&~I3&~I4)|(~I1&I3&I4)|(I0&I3&I4)|(~I0&~I1&~I2&I4)|(~I0&~I1&~I2&I3)|(I0&~I1&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6108  (
            .Z (_N10183_1539),
            .I0 (_N10183_2507),
            .I1 (_N10183_2506),
            .S (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6110  (
            .Z (_N10183_1541),
            .I0 (_N10183_2510),
            .I1 (_N10183_2511),
            .S (\u_lcd_rgb_char/bcd_data_x [13] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6111  (
            .Z (_N10183_1542),
            .I0 (_N10183_2512),
            .I1 (_N10183_2513),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6112  (
            .Z (_N10183_1543),
            .I0 (_N10183_2515),
            .I1 (_N10183_2514),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6113  (
            .Z (_N10183_1544),
            .I0 (_N10183_2517),
            .I1 (_N10183_2516),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6115  */ #(
            .INIT(32'b11111110111110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6115  (
            .Z (_N10183_1546),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (_N10183_2520));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I2&I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6116  */ #(
            .INIT(32'b11101111111111111010101010101010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6116  (
            .Z (_N10183_1547),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .ID (_N10183_2521));
	// LUT = (ID&~I4)|(~I3&I4)|(~I2&I4)|(I1&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6119  */ #(
            .INIT(32'b10111111110110011101101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6119  (
            .Z (_N10183_1550),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&I2&~I4)|(~I2&I3&I4)|(I0&I3&I4)|(~I0&I2&~I3)|(I0&~I2&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6120  */ #(
            .INIT(32'b10011000010110100111010011000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6120  (
            .Z (_N10183_1551),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&I2&~I3&~I4)|(~I1&I2&I3&~I4)|(~I0&I1&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I2&I4)|(I0&~I1&~I2&~I3)|(~I0&I1&I2&~I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6124  */ #(
            .INIT(32'b10111011111100111011101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6124  (
            .Z (_N10183_1555),
            .I0 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(I2&~I3)|(I0&I3)|(~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6126  */ #(
            .INIT(32'b10011111100111101111100111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6126  (
            .Z (_N10183_1557),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2&~I4)|(I1&~I2&I4)|(I0&~I2&I4)|(I1&~I2&~I3)|(I0&~I2&~I3)|(~I0&~I1&I3)|(~I0&~I1&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6129  */ #(
            .INIT(32'b11101000111111101110111111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6129  (
            .Z (_N10183_1560),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (_N10183_3460));
	// LUT = (~I2&~I4)|(ID&~I4)|(I2&~I3&I4)|(I0&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I1&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6130  */ #(
            .INIT(32'b10101010101010101110011001000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6130  (
            .Z (_N10183_1561),
            .I0 (_N10183_2539),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [12] ));
	// LUT = (ID&I2&I3&~I4)|(ID&~I1&I3&~I4)|(~ID&I1&I3&~I4)|(~ID&I1&I2&~I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6132  */ #(
            .INIT(32'b11101100111011001101101110011011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6132  (
            .Z (_N10183_1563),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I2&~I4)|(~I0&~I1&~I4)|(I0&I2&I4)|(I1&I4)|(I1&I2&I3)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6138  */ #(
            .INIT(32'b11110111110001111101001111110011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6138  (
            .Z (_N10183_1569),
            .I0 (_N10183_2712),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .ID (_N10183_2642));
	// LUT = (~I1&~I3&~I4)|(~I1&I3&I4)|(~I0&I1&I4)|(~ID&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6140  */ #(
            .INIT(32'b11001100001100110000110100100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6140  (
            .Z (_N10183_1571),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I2&I3&~I4)|(~I1&~I3&I4)|(I1&I3&I4)|(I0&~I1&I2&~I3)|(I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6141  */ #(
            .INIT(32'b11110110111111101111100010011000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6141  (
            .Z (_N10183_1572),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I4)|(I0&~I1&I4)|(~I0&I1&I4)|(I0&I1&~I3)|(I2&I3)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6143  */ #(
            .INIT(32'b11101111011011110000100101101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6143  (
            .Z (_N10183_1574),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I0&I1&I4)|(I0&~I1&~I3)|(~I0&I1&~I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6145  */ #(
            .INIT(32'b10100101101001010001000100000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6145  (
            .Z (_N10183_1576),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I3&~I4)|(~I0&~I2&I4)|(I0&I2&I4)|(~I0&~I1&~I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6146_3  */ #(
            .INIT(32'b11001100000100011111111111111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6146_3  (
            .Z (_N10183_1577),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (_N10183_1004));
	// LUT = (I3&~I4)|(I2&~I4)|(I1&~I4)|(~ID&~I4)|(~I0&~I1&~I3&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6147  */ #(
            .INIT(32'b11110101000100010100010011110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6147  (
            .Z (_N10183_1578),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = (I2&~I3&~I4)|(~I0&I1&~I4)|(I2&I3&I4)|(~I0&~I1&I4)|(~I0&~I1&~I3)|(~I0&I1&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6150  (
            .Z (_N10183_1581),
            .I0 (_N10183_2569),
            .I1 (_N10183_2570),
            .S (\u_lcd_rgb_char/bcd_data_x [13] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6153  */ #(
            .INIT(32'b11111111101100110101100111101101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6153  (
            .Z (_N10183_1584),
            .I0 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(ID&~I1&I2&~I3)|(I0&ID&I2&~I3)|(ID&I1&~I2&I3)|(~ID&I2&I3)|(~ID&~I1&~I2)|(I0&~ID&I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6154  */ #(
            .INIT(32'b10101010101010101100111011001100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6154  (
            .Z (_N10183_1585),
            .I0 (_N10183_2577),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [13] ));
	// LUT = (ID&~I2&I3&~I4)|(I1&~I4)|(I0&I4) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6156  */ #(
            .INIT(32'b11011110000100101101110000010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6156  (
            .Z (_N10183_1587),
            .I0 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I3 (_N10183_2579),
            .I4 (_N10183_1748),
            .ID (\u_lcd_rgb_char/bcd_data_x [12] ));
	// LUT = (~ID&~I1&I2&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6157  */ #(
            .INIT(32'b10101000011010000000001000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6157  (
            .Z (_N10183_1588),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&I1&I2&~I3&I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(I0&~I1&I2&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6159  */ #(
            .INIT(32'b10100101111100011110001001011010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6159  (
            .Z (_N10183_1590),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I3&~I4)|(I0&~I1&~I2&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I3&I4)|(~I0&~I1&~I2&I4)|(I0&I2&I4)|(~I0&I2&~I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6160  */ #(
            .INIT(32'b11101010110010001100101010010100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6160  (
            .Z (_N10183_1591),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&~I2&~I3&~I4)|(~I0&~I1&I2&~I3&~I4)|(I0&I3&I4)|(I1&I2&I4)|(I0&I1&I4)|(I0&~I2&I3)|(I1&I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6161  */ #(
            .INIT(32'b10100010111100101111111100101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6161  (
            .Z (_N10183_1592),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3&~I4)|(~I2&~I4)|(I2&~I3&I4)|(I0&I2&I3)|(I0&~I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6165  (
            .Z (_N10183_1596),
            .I0 (_N10183_2592),
            .I1 (_N10183_2593),
            .S (\u_lcd_rgb_char/bcd_data_x [15] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6166  (
            .Z (_N10183_1597),
            .I0 (_N10183_2594),
            .I1 (_N10183_2595),
            .S (\u_lcd_rgb_char/bcd_data_x [13] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6167  (
            .Z (_N10183_1598),
            .I0 (_N10183_2597),
            .I1 (_N10183_2596),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6169  */ #(
            .INIT(32'b11110011111011111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6169  (
            .Z (_N10183_1600),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I4)|(~I0&~I4)|(I0&~I1&I4)|(I1&~I3)|(~I0&~I1&I3)|(~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6172  */ #(
            .INIT(32'b10011011000100111001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6172  (
            .Z (_N10183_1603),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I1&~I2&~I4)|(~I1&~I2&I4)|(~I0&~I1&I4)|(~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6173  */ #(
            .INIT(16'b1001100100001001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6173  (
            .Z (_N10183_1604),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3)|(I0&I1&I3)|(~I0&~I1&~I2)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6175  */ #(
            .INIT(32'b11111111110110111101111111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6175  (
            .Z (_N10183_1606),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I4)|(I3&I4)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6176  */ #(
            .INIT(32'b11011111111011111110101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6176  (
            .Z (_N10183_1607),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I4)|(~I0&I3&I4)|(I1&~I3)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6177  */ #(
            .INIT(32'b11111011111011111110011111101011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6177  (
            .Z (_N10183_1608),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&I3&~I4)|(I1&~I3&I4)|(~I1&I3&I4)|(I0&I4)|(I0&~I3)|(~I1&~I2)|(I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6179  */ #(
            .INIT(32'b11111000000000000001111000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6179  (
            .Z (_N10183_1610),
            .I0 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&~I2&I3&~I4)|(I0&~I2&~I4)|(I2&I3&I4)|(I0&I1&~I2&I3)|(~I0&~I1&I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6181  */ #(
            .INIT(32'b10101000101010000101001000001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6181  (
            .Z (_N10183_1612),
            .I0 (_N10183_3516),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .ID (\u_lcd_rgb_char/bcd_data_x [14] ));
	// LUT = (ID&~I2&~I3&~I4)|(~ID&I2&I3&~I4)|(ID&~I1&~I2&~I4)|(I0&I2&I4)|(I0&I1&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_6182  (
            .Z (_N10183_1613),
            .I0 (_N10183_2621),
            .I1 (_N10183_2620),
            .S (\u_lcd_rgb_char/pixel_xpos_w [2] ));

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_6184  */ #(
            .INIT(32'b10101011101110110101010101010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6184  (
            .Z (_N10183_1615),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .ID (_N10183_2623));
	// LUT = (~ID&~I4)|(~I1&~I3&I4)|(~I1&~I2&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6191  */ #(
            .INIT(32'b11100000000000000110001000010001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6191  (
            .Z (_N10183_1622),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I0&~I1&I3&~I4)|(I0&I2&I3&I4)|(~I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6192  */ #(
            .INIT(32'b10010001011101111110111100010111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6192  (
            .Z (_N10183_1623),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&I3&~I4)|(I0&I3&~I4)|(~I1&~I3&I4)|(~I0&~I3&I4)|(~I0&~I1&I4)|(~I1&~I2&~I3)|(~I0&~I2&~I3)|(~I0&~I1&~I3)|(I0&I1&I2&I3)|(~I0&~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6194  */ #(
            .INIT(32'b11111111001000000011111110100000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6194  (
            .Z (_N10183_1625),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I0&I2&~I3&~I4)|(I3&I4)|(~I2&I3)|(~I1&I3)|(I0&~I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_6203  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6203  (
            .Z (_N10183_1634),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = I0&I1 ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6225  */ #(
            .INIT(16'b1010100001000100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6225  (
            .Z (_N10183_1656),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I1&~I3)|(I0&I2&I3)|(I0&I1&I3) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_6226  */ #(
            .INIT(8'b11101000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6226  (
            .Z (_N10183_1657),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&I2)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6237  */ #(
            .INIT(32'b11101101111111011010110001010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6237  (
            .Z (_N10183_1668),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(I0&I2&I3)|(I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6240  */ #(
            .INIT(32'b11101101010101011010101110111001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6240  (
            .Z (_N10183_1671),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I3&~I4)|(I0&I2&~I4)|(I0&I1&~I4)|(~I0&I1&I4)|(~I0&~I1&~I3)|(I0&I2&I3)|(I0&I1&I3)|(~I0&~I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6241  */ #(
            .INIT(32'b11111101111111111110111110111001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6241  (
            .Z (_N10183_1672),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I3&~I4)|(~I3&I4)|(~I0&I4)|(~I0&~I1&~I3)|(I1&I3)|(~I0&~I1&~I2)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6242  */ #(
            .INIT(32'b10111010001000100100011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6242  (
            .Z (_N10183_1673),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I2&~I3&~I4)|(~I0&I1&I3&~I4)|(~I1&I2&I3&I4)|(I0&I3&I4)|(I0&~I1&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6243  */ #(
            .INIT(32'b11111111111101111110111111011110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6243  (
            .Z (_N10183_1674),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(~I1&I4)|(~I0&I2&~I3)|(~I2&I3)|(I0&I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6245  */ #(
            .INIT(32'b11100101111111111011101011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6245  (
            .Z (_N10183_1676),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I1&I2&I3&~I4)|(I0&~I4)|(~I3&I4)|(~I0&~I2&I4)|(~I0&I1&I4)|(I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6246  */ #(
            .INIT(32'b10111001110111101111111111001110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6246  (
            .Z (_N10183_1677),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I4)|(I1&~I4)|(~I0&~I1&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I0&I2&I3)|(~I0&~I1&I3)|(I0&I1) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6247_5  */ #(
            .INIT(16'b1111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6247_5  (
            .Z (_N10183_1678),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6249  */ #(
            .INIT(32'b10011010100100111110101111101001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6249  (
            .Z (_N10183_1680),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I2&~I4)|(I1&I2&~I4)|(I0&I2&~I4)|(I0&I1&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(~I0&~I1&~I2&~I3)|(I0&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6250  */ #(
            .INIT(32'b11111101111011110000011010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6250  (
            .Z (_N10183_1681),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(I0&~I3&I4)|(~I0&I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6251  */ #(
            .INIT(32'b11110111111111010000010010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6251  (
            .Z (_N10183_1682),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&I4)|(~I1&I3&I4)|(I2&I4)|(~I0&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6254  */ #(
            .INIT(32'b11001001110001000000001100001101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6254  (
            .Z (_N10183_1685),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(~I0&~I1&~I2&~I4)|(I0&I1&I3&I4)|(I1&I2&I4)|(~I0&I1&~I2&~I3)|(~I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6275  */ #(
            .INIT(32'b11001100000000010001011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6275  (
            .Z (_N10183_1706),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&~I1&I2&I3&~I4)|(I1&I3&I4)|(~I0&~I1&~I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6276  */ #(
            .INIT(16'b1101100001001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6276  (
            .Z (_N10183_1707),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&I2&I3)|(I0&I1&I3)|(I0&I1&~I2)|(~I0&I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_6285  */ #(
            .INIT(4'b1001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6285  (
            .Z (_N10183_1716),
            .I0 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = ~I1^I0 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6308  */ #(
            .INIT(32'b11011111101010111111111010111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6308  (
            .Z (_N10183_1739),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I2&~I4)|(~I1&I2&~I4)|(~I1&~I2&I4)|(~I1&~I2&~I3)|(I0&~I3)|(~I0&I2&I3)|(I1&I3)|(I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6309  */ #(
            .INIT(32'b11111111010111101110010010101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6309  (
            .Z (_N10183_1740),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I2&~I4)|(I3&I4)|(~I0&I2&I4)|(I0&~I2&~I3)|(~I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6310  */ #(
            .INIT(32'b11110010000000001000101100010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6310  (
            .Z (_N10183_1741),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(I0&I1&I3&~I4)|(I2&I3&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6311  */ #(
            .INIT(32'b10010000011001101001000101100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6311  (
            .Z (_N10183_1742),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3&~I4)|(I0&~I1&~I3&I4)|(I0&~I1&I2&~I3)|(~I0&I1&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6316  */ #(
            .INIT(32'b11111111110111111111101111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6316  (
            .Z (_N10183_1747),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_6317  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6317  (
            .Z (_N10183_1748),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6318  */ #(
            .INIT(32'b11111110111111111101011011110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6318  (
            .Z (_N10183_1749),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I4)|(~I1&~I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6319  */ #(
            .INIT(32'b10111001000111010111100001000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6319  (
            .Z (_N10183_1750),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I4)|(~I0&I1&~I2&~I3)|(I0&I1&~I2&I3)|(~I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6333  */ #(
            .INIT(32'b11001100111111101010111010100011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6333  (
            .Z (_N10183_1764),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&~I2&~I3&~I4)|(I0&~I1&~I4)|(I2&~I3&I4)|(I1&I4)|(I0&~I1&~I3)|(I1&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6334  */ #(
            .INIT(32'b11110010001100111111101111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6334  (
            .Z (_N10183_1765),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I3&~I4)|(~I1&I3&~I4)|(I0&~I4)|(~I1&~I3&I4)|(I2&I3)|(~I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6335  */ #(
            .INIT(32'b11111110111111101110111000010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6335  (
            .Z (_N10183_1766),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I2&I4)|(I0&I4)|(I1&I3)|(I0&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6336  */ #(
            .INIT(32'b10110011001101111111101100001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6336  (
            .Z (_N10183_1767),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&~I2&~I4)|(~I0&~I2&~I3&I4)|(~I1&I4)|(I0&I2&I3)|(~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6337  */ #(
            .INIT(32'b11111011111111111111101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6337  (
            .Z (_N10183_1768),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I3&I4)|(I2)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6338  */ #(
            .INIT(32'b10111011101110111111101110011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6338  (
            .Z (_N10183_1769),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&I4)|(I0&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6360  */ #(
            .INIT(32'b11111100111111111100000011110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6360  (
            .Z (_N10183_1791),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I4)|(I1&I4)|(~I1&~I3)|(~I0&~I3)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6365  */ #(
            .INIT(32'b10111111101111111101010101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6365  (
            .Z (_N10183_1796),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I4)|(I0&I4)|(~I2&~I3)|(I0&I1&I2&I3)|(~I0&~I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6368  */ #(
            .INIT(32'b10100101101001010100000001001111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6368  (
            .Z (_N10183_1799),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I4)|(I0&I2&I4) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6372  */ #(
            .INIT(16'b1100100110010011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6372  (
            .Z (_N10183_1803),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I1&~I2&~I3)|(~I0&~I1&~I3)|(I1&I2&I3)|(I0&I1&I3)|(~I0&~I1&~I2)|(I0&I1&I2) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6374  */ #(
            .INIT(16'b1011111110110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6374  (
            .Z (_N10183_1805),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3)|(~I0&~I2)|(I0&I2)|(~I0&~I1) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_6375  */ #(
            .INIT(8'b11001101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6375  (
            .Z (_N10183_1806),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (~I0&~I2)|(I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6387  */ #(
            .INIT(32'b11101101111111011010110001010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6387  (
            .Z (_N10183_1818),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(I0&I2&I3)|(I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6390  */ #(
            .INIT(32'b11101101111111010101010111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6390  (
            .Z (_N10183_1821),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&~I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(~I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6391  */ #(
            .INIT(32'b10101011111011111011100110111001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6391  (
            .Z (_N10183_1822),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I4)|(I1&~I3&I4)|(I0&I4)|(~I0&~I1&~I2)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6392  */ #(
            .INIT(32'b10111010001000100100011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6392  (
            .Z (_N10183_1823),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I2&~I3&~I4)|(~I0&I1&I3&~I4)|(~I1&I2&I3&I4)|(I0&I3&I4)|(I0&~I1&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6393  */ #(
            .INIT(32'b11111111111101111110111111011110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6393  (
            .Z (_N10183_1824),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(~I1&I4)|(~I0&I2&~I3)|(~I2&I3)|(I0&I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6395  */ #(
            .INIT(32'b11100101111111111011101011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6395  (
            .Z (_N10183_1826),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I1&I2&I3&~I4)|(I0&~I4)|(~I3&I4)|(~I0&~I2&I4)|(~I0&I1&I4)|(I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6396  */ #(
            .INIT(32'b10111001110111101111111111001110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6396  (
            .Z (_N10183_1827),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I4)|(I1&~I4)|(~I0&~I1&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I0&I2&I3)|(~I0&~I1&I3)|(I0&I1) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6397_3  */ #(
            .INIT(16'b1111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6397_3  (
            .Z (_N10183_1828),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6399  */ #(
            .INIT(32'b10011010100100111110101111101001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6399  (
            .Z (_N10183_1830),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I2&~I4)|(I1&I2&~I4)|(I0&I2&~I4)|(I0&I1&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(~I0&~I1&~I2&~I3)|(I0&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6400  */ #(
            .INIT(32'b11111101111011110000011010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6400  (
            .Z (_N10183_1831),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(I0&~I3&I4)|(~I0&I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6401  */ #(
            .INIT(32'b11110111111111010000010010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6401  (
            .Z (_N10183_1832),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&I4)|(~I1&I3&I4)|(I2&I4)|(~I0&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6404  */ #(
            .INIT(32'b11001001110001000000001100001101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6404  (
            .Z (_N10183_1835),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(~I0&~I1&~I2&~I4)|(I0&I1&I3&I4)|(I1&I2&I4)|(~I0&I1&~I2&~I3)|(~I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6423  */ #(
            .INIT(32'b11001100000000010001011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6423  (
            .Z (_N10183_1854),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&~I1&I2&I3&~I4)|(I1&I3&I4)|(~I0&~I1&~I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6424  */ #(
            .INIT(16'b1101100001001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6424  (
            .Z (_N10183_1855),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&I2&I3)|(I0&I1&I3)|(I0&I1&~I2)|(~I0&I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_6432  */ #(
            .INIT(4'b1001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6432  (
            .Z (_N10183_1863),
            .I0 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = ~I1^I0 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6453  */ #(
            .INIT(32'b11011111101010111111111010111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6453  (
            .Z (_N10183_1884),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I2&~I4)|(~I1&I2&~I4)|(~I1&~I2&I4)|(~I1&~I2&~I3)|(I0&~I3)|(~I0&I2&I3)|(I1&I3)|(I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6454  */ #(
            .INIT(32'b11111111010111101110010010101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6454  (
            .Z (_N10183_1885),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I2&~I4)|(I3&I4)|(~I0&I2&I4)|(I0&~I2&~I3)|(~I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6455  */ #(
            .INIT(32'b11110010000000001000101100010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6455  (
            .Z (_N10183_1886),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(I0&I1&I3&~I4)|(I2&I3&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6456  */ #(
            .INIT(32'b10010000011001101001000101100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6456  (
            .Z (_N10183_1887),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3&~I4)|(I0&~I1&~I3&I4)|(I0&~I1&I2&~I3)|(~I0&I1&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6461  */ #(
            .INIT(32'b11111111110111111111101111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6461  (
            .Z (_N10183_1892),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6462  */ #(
            .INIT(32'b11111110111111111101011011110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6462  (
            .Z (_N10183_1893),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I4)|(~I1&~I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6463  */ #(
            .INIT(32'b10111001000111010111100001000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6463  (
            .Z (_N10183_1894),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I4)|(~I0&I1&~I2&~I3)|(I0&I1&~I2&I3)|(~I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6476  */ #(
            .INIT(32'b11001100111111101010111010100011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6476  (
            .Z (_N10183_1907),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&~I2&~I3&~I4)|(I0&~I1&~I4)|(I2&~I3&I4)|(I1&I4)|(I0&~I1&~I3)|(I1&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6477  */ #(
            .INIT(32'b11110010001100111111101111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6477  (
            .Z (_N10183_1908),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I3&~I4)|(~I1&I3&~I4)|(I0&~I4)|(~I1&~I3&I4)|(I2&I3)|(~I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6478  */ #(
            .INIT(32'b11111110111111101110111000010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6478  (
            .Z (_N10183_1909),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I2&I4)|(I0&I4)|(I1&I3)|(I0&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6479  */ #(
            .INIT(32'b10110011001101111111101100001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6479  (
            .Z (_N10183_1910),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&~I2&~I4)|(~I0&~I2&~I3&I4)|(~I1&I4)|(I0&I2&I3)|(~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6480  */ #(
            .INIT(32'b11111011111111111111101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6480  (
            .Z (_N10183_1911),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I3&I4)|(I2)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6481  */ #(
            .INIT(32'b10111011101110111111101110011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6481  (
            .Z (_N10183_1912),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&I4)|(I0&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6505  */ #(
            .INIT(32'b10111111101111111101010101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6505  (
            .Z (_N10183_1936),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I4)|(I0&I4)|(~I2&~I3)|(I0&I1&I2&I3)|(~I0&~I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6507  */ #(
            .INIT(32'b10100101101001010100000001001111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6507  (
            .Z (_N10183_1938),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I4)|(I0&I2&I4) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6512  */ #(
            .INIT(16'b1011111110110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6512  (
            .Z (_N10183_1943),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3)|(~I0&~I2)|(I0&I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6524  */ #(
            .INIT(32'b11101101111111011010110001010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6524  (
            .Z (_N10183_1955),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(I0&I2&I3)|(I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6527  */ #(
            .INIT(32'b11101101111111010101010111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6527  (
            .Z (_N10183_1958),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&~I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(~I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6528  */ #(
            .INIT(32'b10101011111011111011100110111001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6528  (
            .Z (_N10183_1959),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I4)|(I1&~I3&I4)|(I0&I4)|(~I0&~I1&~I2)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6529  */ #(
            .INIT(32'b10111010001000100100011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6529  (
            .Z (_N10183_1960),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I2&~I3&~I4)|(~I0&I1&I3&~I4)|(~I1&I2&I3&I4)|(I0&I3&I4)|(I0&~I1&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6530  */ #(
            .INIT(32'b11111111111101111110111111011110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6530  (
            .Z (_N10183_1961),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(~I1&I4)|(~I0&I2&~I3)|(~I2&I3)|(I0&I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6532  */ #(
            .INIT(32'b11100101111111111011101011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6532  (
            .Z (_N10183_1963),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I1&I2&I3&~I4)|(I0&~I4)|(~I3&I4)|(~I0&~I2&I4)|(~I0&I1&I4)|(I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6533  */ #(
            .INIT(32'b10111001110111101111111111001110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6533  (
            .Z (_N10183_1964),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I4)|(I1&~I4)|(~I0&~I1&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I0&I2&I3)|(~I0&~I1&I3)|(I0&I1) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6534_3  */ #(
            .INIT(16'b1111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6534_3  (
            .Z (_N10183_1965),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6536  */ #(
            .INIT(32'b10011010100100111110101111101001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6536  (
            .Z (_N10183_1967),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I2&~I4)|(I1&I2&~I4)|(I0&I2&~I4)|(I0&I1&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(~I0&~I1&~I2&~I3)|(I0&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6537  */ #(
            .INIT(32'b11111101111011110000011010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6537  (
            .Z (_N10183_1968),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(I0&~I3&I4)|(~I0&I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6538  */ #(
            .INIT(32'b11110111111111010000010010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6538  (
            .Z (_N10183_1969),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&I4)|(~I1&I3&I4)|(I2&I4)|(~I0&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6541  */ #(
            .INIT(32'b11001001110001000000001100001101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6541  (
            .Z (_N10183_1972),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(~I0&~I1&~I2&~I4)|(I0&I1&I3&I4)|(I1&I2&I4)|(~I0&I1&~I2&~I3)|(~I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6560  */ #(
            .INIT(32'b11001100000000010001011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6560  (
            .Z (_N10183_1991),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&~I1&I2&I3&~I4)|(I1&I3&I4)|(~I0&~I1&~I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6561  */ #(
            .INIT(16'b1101100001001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6561  (
            .Z (_N10183_1992),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&I2&I3)|(I0&I1&I3)|(I0&I1&~I2)|(~I0&I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_6569  */ #(
            .INIT(4'b1001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6569  (
            .Z (_N10183_2000),
            .I0 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = ~I1^I0 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6590  */ #(
            .INIT(32'b11011111101010111111111010111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6590  (
            .Z (_N10183_2021),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I2&~I4)|(~I1&I2&~I4)|(~I1&~I2&I4)|(~I1&~I2&~I3)|(I0&~I3)|(~I0&I2&I3)|(I1&I3)|(I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6591  */ #(
            .INIT(32'b11111111010111101110010010101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6591  (
            .Z (_N10183_2022),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I2&~I4)|(I3&I4)|(~I0&I2&I4)|(I0&~I2&~I3)|(~I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6592  */ #(
            .INIT(32'b11110010000000001000101100010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6592  (
            .Z (_N10183_2023),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(I0&I1&I3&~I4)|(I2&I3&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6593  */ #(
            .INIT(32'b10010000011001101001000101100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6593  (
            .Z (_N10183_2024),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3&~I4)|(I0&~I1&~I3&I4)|(I0&~I1&I2&~I3)|(~I0&I1&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6598  */ #(
            .INIT(32'b11111111110111111111101111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6598  (
            .Z (_N10183_2029),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6599  */ #(
            .INIT(32'b11111110111111111101011011110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6599  (
            .Z (_N10183_2030),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I4)|(~I1&~I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6600  */ #(
            .INIT(32'b10111001000111010111100001000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6600  (
            .Z (_N10183_2031),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I4)|(~I0&I1&~I2&~I3)|(I0&I1&~I2&I3)|(~I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6613  */ #(
            .INIT(32'b11001100111111101010111010100011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6613  (
            .Z (_N10183_2044),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&~I2&~I3&~I4)|(I0&~I1&~I4)|(I2&~I3&I4)|(I1&I4)|(I0&~I1&~I3)|(I1&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6614  */ #(
            .INIT(32'b11110010001100111111101111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6614  (
            .Z (_N10183_2045),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I3&~I4)|(~I1&I3&~I4)|(I0&~I4)|(~I1&~I3&I4)|(I2&I3)|(~I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6615  */ #(
            .INIT(32'b11111110111111101110111000010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6615  (
            .Z (_N10183_2046),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I2&I4)|(I0&I4)|(I1&I3)|(I0&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6616  */ #(
            .INIT(32'b10110011001101111111101100001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6616  (
            .Z (_N10183_2047),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&~I2&~I4)|(~I0&~I2&~I3&I4)|(~I1&I4)|(I0&I2&I3)|(~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6617  */ #(
            .INIT(32'b11111011111111111111101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6617  (
            .Z (_N10183_2048),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I3&I4)|(I2)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6618  */ #(
            .INIT(32'b10111011101110111111101110011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6618  (
            .Z (_N10183_2049),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&I4)|(I0&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6642  */ #(
            .INIT(32'b10111111101111111101010101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6642  (
            .Z (_N10183_2073),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I4)|(I0&I4)|(~I2&~I3)|(I0&I1&I2&I3)|(~I0&~I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6644  */ #(
            .INIT(32'b10100101101001010100000001001111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6644  (
            .Z (_N10183_2075),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I4)|(I0&I2&I4) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6649  */ #(
            .INIT(16'b1011111110110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6649  (
            .Z (_N10183_2080),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3)|(~I0&~I2)|(I0&I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6661  */ #(
            .INIT(32'b11101101111111011010110001010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6661  (
            .Z (_N10183_2092),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(I0&I2&I3)|(I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6664  */ #(
            .INIT(32'b11101101111111010101010111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6664  (
            .Z (_N10183_2095),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&~I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(~I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6665  */ #(
            .INIT(32'b10101011111011111011100110111001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6665  (
            .Z (_N10183_2096),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I4)|(I1&~I3&I4)|(I0&I4)|(~I0&~I1&~I2)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6666  */ #(
            .INIT(32'b10111010001000100100011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6666  (
            .Z (_N10183_2097),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I2&~I3&~I4)|(~I0&I1&I3&~I4)|(~I1&I2&I3&I4)|(I0&I3&I4)|(I0&~I1&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6667  */ #(
            .INIT(32'b11111111111101111110111111011110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6667  (
            .Z (_N10183_2098),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(~I1&I4)|(~I0&I2&~I3)|(~I2&I3)|(I0&I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6669  */ #(
            .INIT(32'b11100101111111111011101011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6669  (
            .Z (_N10183_2100),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I1&I2&I3&~I4)|(I0&~I4)|(~I3&I4)|(~I0&~I2&I4)|(~I0&I1&I4)|(I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6670  */ #(
            .INIT(32'b10111001110111101111111111001110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6670  (
            .Z (_N10183_2101),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I4)|(I1&~I4)|(~I0&~I1&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I0&I2&I3)|(~I0&~I1&I3)|(I0&I1) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6671_3  */ #(
            .INIT(16'b1111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6671_3  (
            .Z (_N10183_2102),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6673  */ #(
            .INIT(32'b10011010100100111110101111101001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6673  (
            .Z (_N10183_2104),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I2&~I4)|(I1&I2&~I4)|(I0&I2&~I4)|(I0&I1&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(~I0&~I1&~I2&~I3)|(I0&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6674  */ #(
            .INIT(32'b11111101111011110000011010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6674  (
            .Z (_N10183_2105),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(I0&~I3&I4)|(~I0&I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6675  */ #(
            .INIT(32'b11110111111111010000010010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6675  (
            .Z (_N10183_2106),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&I4)|(~I1&I3&I4)|(I2&I4)|(~I0&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6678  */ #(
            .INIT(32'b11001001110001000000001100001101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6678  (
            .Z (_N10183_2109),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(~I0&~I1&~I2&~I4)|(I0&I1&I3&I4)|(I1&I2&I4)|(~I0&I1&~I2&~I3)|(~I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6697  */ #(
            .INIT(32'b11001100000000010001011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6697  (
            .Z (_N10183_2128),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&~I1&I2&I3&~I4)|(I1&I3&I4)|(~I0&~I1&~I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6698  */ #(
            .INIT(16'b1101100001001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6698  (
            .Z (_N10183_2129),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&I2&I3)|(I0&I1&I3)|(I0&I1&~I2)|(~I0&I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_6706  */ #(
            .INIT(4'b1001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6706  (
            .Z (_N10183_2137),
            .I0 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = ~I1^I0 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6727  */ #(
            .INIT(32'b11011111101010111111111010111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6727  (
            .Z (_N10183_2158),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I2&~I4)|(~I1&I2&~I4)|(~I1&~I2&I4)|(~I1&~I2&~I3)|(I0&~I3)|(~I0&I2&I3)|(I1&I3)|(I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6728  */ #(
            .INIT(32'b11111111010111101110010010101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6728  (
            .Z (_N10183_2159),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I2&~I4)|(I3&I4)|(~I0&I2&I4)|(I0&~I2&~I3)|(~I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6729  */ #(
            .INIT(32'b11110010000000001000101100010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6729  (
            .Z (_N10183_2160),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(I0&I1&I3&~I4)|(I2&I3&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6730  */ #(
            .INIT(32'b10010000011001101001000101100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6730  (
            .Z (_N10183_2161),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3&~I4)|(I0&~I1&~I3&I4)|(I0&~I1&I2&~I3)|(~I0&I1&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6735  */ #(
            .INIT(32'b11111111110111111111101111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6735  (
            .Z (_N10183_2166),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6736  */ #(
            .INIT(32'b11111110111111111101011011110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6736  (
            .Z (_N10183_2167),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I4)|(~I1&~I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6737  */ #(
            .INIT(32'b10111001000111010111100001000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6737  (
            .Z (_N10183_2168),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I4)|(~I0&I1&~I2&~I3)|(I0&I1&~I2&I3)|(~I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6750  */ #(
            .INIT(32'b11001100111111101010111010100011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6750  (
            .Z (_N10183_2181),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&~I2&~I3&~I4)|(I0&~I1&~I4)|(I2&~I3&I4)|(I1&I4)|(I0&~I1&~I3)|(I1&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6751  */ #(
            .INIT(32'b11110010001100111111101111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6751  (
            .Z (_N10183_2182),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I3&~I4)|(~I1&I3&~I4)|(I0&~I4)|(~I1&~I3&I4)|(I2&I3)|(~I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6752  */ #(
            .INIT(32'b11111110111111101110111000010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6752  (
            .Z (_N10183_2183),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I2&I4)|(I0&I4)|(I1&I3)|(I0&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6753  */ #(
            .INIT(32'b10110011001101111111101100001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6753  (
            .Z (_N10183_2184),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&~I2&~I4)|(~I0&~I2&~I3&I4)|(~I1&I4)|(I0&I2&I3)|(~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6754  */ #(
            .INIT(32'b11111011111111111111101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6754  (
            .Z (_N10183_2185),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I3&I4)|(I2)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6755  */ #(
            .INIT(32'b10111011101110111111101110011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6755  (
            .Z (_N10183_2186),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&I4)|(I0&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6779  */ #(
            .INIT(32'b10111111101111111101010101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6779  (
            .Z (_N10183_2210),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I4)|(I0&I4)|(~I2&~I3)|(I0&I1&I2&I3)|(~I0&~I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6781  */ #(
            .INIT(32'b10100101101001010100000001001111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6781  (
            .Z (_N10183_2212),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I4)|(I0&I2&I4) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6786  */ #(
            .INIT(16'b1011111110110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6786  (
            .Z (_N10183_2217),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3)|(~I0&~I2)|(I0&I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6798  */ #(
            .INIT(32'b11101101111111011010110001010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6798  (
            .Z (_N10183_2229),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(I0&I2&I3)|(I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6801  */ #(
            .INIT(32'b11101101111111010101010111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6801  (
            .Z (_N10183_2232),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&~I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(~I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6802  */ #(
            .INIT(32'b10101011111011111011100110111001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6802  (
            .Z (_N10183_2233),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I4)|(I1&~I3&I4)|(I0&I4)|(~I0&~I1&~I2)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6803  */ #(
            .INIT(32'b10111010001000100100011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6803  (
            .Z (_N10183_2234),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I2&~I3&~I4)|(~I0&I1&I3&~I4)|(~I1&I2&I3&I4)|(I0&I3&I4)|(I0&~I1&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6804  */ #(
            .INIT(32'b11111111111101111110111111011110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6804  (
            .Z (_N10183_2235),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(~I1&I4)|(~I0&I2&~I3)|(~I2&I3)|(I0&I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6806  */ #(
            .INIT(32'b11100101111111111011101011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6806  (
            .Z (_N10183_2237),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I1&I2&I3&~I4)|(I0&~I4)|(~I3&I4)|(~I0&~I2&I4)|(~I0&I1&I4)|(I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6807  */ #(
            .INIT(32'b10111001110111101111111111001110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6807  (
            .Z (_N10183_2238),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I4)|(I1&~I4)|(~I0&~I1&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I0&I2&I3)|(~I0&~I1&I3)|(I0&I1) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6808_3  */ #(
            .INIT(16'b1111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6808_3  (
            .Z (_N10183_2239),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6810  */ #(
            .INIT(32'b10011010100100111110101111101001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6810  (
            .Z (_N10183_2241),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I2&~I4)|(I1&I2&~I4)|(I0&I2&~I4)|(I0&I1&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(~I0&~I1&~I2&~I3)|(I0&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6811  */ #(
            .INIT(32'b11111101111011110000011010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6811  (
            .Z (_N10183_2242),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(I0&~I3&I4)|(~I0&I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6812  */ #(
            .INIT(32'b11110111111111010000010010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6812  (
            .Z (_N10183_2243),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&I4)|(~I1&I3&I4)|(I2&I4)|(~I0&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6815  */ #(
            .INIT(32'b11001001110001000000001100001101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6815  (
            .Z (_N10183_2246),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(~I0&~I1&~I2&~I4)|(I0&I1&I3&I4)|(I1&I2&I4)|(~I0&I1&~I2&~I3)|(~I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6834  */ #(
            .INIT(32'b11001100000000010001011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6834  (
            .Z (_N10183_2265),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&~I1&I2&I3&~I4)|(I1&I3&I4)|(~I0&~I1&~I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6835  */ #(
            .INIT(16'b1101100001001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6835  (
            .Z (_N10183_2266),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&I2&I3)|(I0&I1&I3)|(I0&I1&~I2)|(~I0&I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_6843  */ #(
            .INIT(4'b1001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6843  (
            .Z (_N10183_2274),
            .I0 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = ~I1^I0 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6864  */ #(
            .INIT(32'b11011111101010111111111010111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6864  (
            .Z (_N10183_2295),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I2&~I4)|(~I1&I2&~I4)|(~I1&~I2&I4)|(~I1&~I2&~I3)|(I0&~I3)|(~I0&I2&I3)|(I1&I3)|(I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6865  */ #(
            .INIT(32'b11111111010111101110010010101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6865  (
            .Z (_N10183_2296),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I2&~I4)|(I3&I4)|(~I0&I2&I4)|(I0&~I2&~I3)|(~I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6866  */ #(
            .INIT(32'b11110010000000001000101100010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6866  (
            .Z (_N10183_2297),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(I0&I1&I3&~I4)|(I2&I3&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6867  */ #(
            .INIT(32'b10010000011001101001000101100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_6867  (
            .Z (_N10183_2298),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3&~I4)|(I0&~I1&~I3&I4)|(I0&~I1&I2&~I3)|(~I0&I1&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6872  */ #(
            .INIT(32'b11111111110111111111101111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6872  (
            .Z (_N10183_2303),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6873  */ #(
            .INIT(32'b11111110111111111101011011110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6873  (
            .Z (_N10183_2304),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I4)|(~I1&~I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6874  */ #(
            .INIT(32'b10111001000111010111100001000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6874  (
            .Z (_N10183_2305),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I4)|(~I0&I1&~I2&~I3)|(I0&I1&~I2&I3)|(~I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6887  */ #(
            .INIT(32'b11001100111111101010111010100011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6887  (
            .Z (_N10183_2318),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&~I2&~I3&~I4)|(I0&~I1&~I4)|(I2&~I3&I4)|(I1&I4)|(I0&~I1&~I3)|(I1&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6888  */ #(
            .INIT(32'b11110010001100111111101111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6888  (
            .Z (_N10183_2319),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I3&~I4)|(~I1&I3&~I4)|(I0&~I4)|(~I1&~I3&I4)|(I2&I3)|(~I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6889  */ #(
            .INIT(32'b11111110111111101110111000010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6889  (
            .Z (_N10183_2320),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I2&I4)|(I0&I4)|(I1&I3)|(I0&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6890  */ #(
            .INIT(32'b10110011001101111111101100001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_6890  (
            .Z (_N10183_2321),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&~I2&~I4)|(~I0&~I2&~I3&I4)|(~I1&I4)|(I0&I2&I3)|(~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6891  */ #(
            .INIT(32'b11111011111111111111101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_6891  (
            .Z (_N10183_2322),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I3&I4)|(I2)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6892  */ #(
            .INIT(32'b10111011101110111111101110011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6892  (
            .Z (_N10183_2323),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&I4)|(I0&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6916  */ #(
            .INIT(32'b10111111101111111101010101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6916  (
            .Z (_N10183_2347),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I4)|(I0&I4)|(~I2&~I3)|(I0&I1&I2&I3)|(~I0&~I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6918  */ #(
            .INIT(32'b10100101101001010100000001001111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6918  (
            .Z (_N10183_2349),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I4)|(I0&I2&I4) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6923  */ #(
            .INIT(16'b1011111110110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6923  (
            .Z (_N10183_2354),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3)|(~I0&~I2)|(I0&I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6935  */ #(
            .INIT(32'b11101101111111011010110001010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6935  (
            .Z (_N10183_2366),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(I0&I2&I3)|(I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6938  */ #(
            .INIT(32'b11101101111111010101010111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_6938  (
            .Z (_N10183_2369),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&~I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(~I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6939  */ #(
            .INIT(32'b10101011111011111011100110111001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6939  (
            .Z (_N10183_2370),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I4)|(I1&~I3&I4)|(I0&I4)|(~I0&~I1&~I2)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6940  */ #(
            .INIT(32'b10111010001000100100011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6940  (
            .Z (_N10183_2371),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I2&~I3&~I4)|(~I0&I1&I3&~I4)|(~I1&I2&I3&I4)|(I0&I3&I4)|(I0&~I1&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6941  */ #(
            .INIT(32'b11111111111101111110111111011110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6941  (
            .Z (_N10183_2372),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(~I1&I4)|(~I0&I2&~I3)|(~I2&I3)|(I0&I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6943  */ #(
            .INIT(32'b11100101111111111011101011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6943  (
            .Z (_N10183_2374),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I1&I2&I3&~I4)|(I0&~I4)|(~I3&I4)|(~I0&~I2&I4)|(~I0&I1&I4)|(I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6944  */ #(
            .INIT(32'b10111001110111101111111111001110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6944  (
            .Z (_N10183_2375),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I4)|(I1&~I4)|(~I0&~I1&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I0&I2&I3)|(~I0&~I1&I3)|(I0&I1) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6945_3  */ #(
            .INIT(16'b1111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_6945_3  (
            .Z (_N10183_2376),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6947  */ #(
            .INIT(32'b10011010100100111110101111101001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6947  (
            .Z (_N10183_2378),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I2&~I4)|(I1&I2&~I4)|(I0&I2&~I4)|(I0&I1&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(~I0&~I1&~I2&~I3)|(I0&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6948  */ #(
            .INIT(32'b11111101111011110000011010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6948  (
            .Z (_N10183_2379),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(I0&~I3&I4)|(~I0&I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6949  */ #(
            .INIT(32'b11110111111111010000010010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6949  (
            .Z (_N10183_2380),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&I4)|(~I1&I3&I4)|(I2&I4)|(~I0&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6952  */ #(
            .INIT(32'b11001001110001000000001100001101))
        \u_lcd_rgb_char/u_lcd_display/N9971_6952  (
            .Z (_N10183_2383),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(~I0&~I1&~I2&~I4)|(I0&I1&I3&I4)|(I1&I2&I4)|(~I0&I1&~I2&~I3)|(~I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_6971  */ #(
            .INIT(32'b11001100000000010001011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6971  (
            .Z (_N10183_2402),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&~I1&I2&I3&~I4)|(I1&I3&I4)|(~I0&~I1&~I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_6972  */ #(
            .INIT(16'b1101100001001000))
        \u_lcd_rgb_char/u_lcd_display/N9971_6972  (
            .Z (_N10183_2403),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&I2&I3)|(I0&I1&I3)|(I0&I1&~I2)|(~I0&I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_6980  */ #(
            .INIT(4'b1001))
        \u_lcd_rgb_char/u_lcd_display/N9971_6980  (
            .Z (_N10183_2411),
            .I0 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = ~I1^I0 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7001  */ #(
            .INIT(32'b11011111101010111111111010111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7001  (
            .Z (_N10183_2432),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I2&~I4)|(~I1&I2&~I4)|(~I1&~I2&I4)|(~I1&~I2&~I3)|(I0&~I3)|(~I0&I2&I3)|(I1&I3)|(I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7002  */ #(
            .INIT(32'b11111111010111101110010010101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7002  (
            .Z (_N10183_2433),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I2&~I4)|(I3&I4)|(~I0&I2&I4)|(I0&~I2&~I3)|(~I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7003  */ #(
            .INIT(32'b11110010000000001000101100010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_7003  (
            .Z (_N10183_2434),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(I0&I1&I3&~I4)|(I2&I3&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7004  */ #(
            .INIT(32'b10010000011001101001000101100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_7004  (
            .Z (_N10183_2435),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3&~I4)|(I0&~I1&~I3&I4)|(I0&~I1&I2&~I3)|(~I0&I1&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7009  */ #(
            .INIT(32'b11111111110111111111101111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7009  (
            .Z (_N10183_2440),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7010  */ #(
            .INIT(32'b11111110111111111101011011110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7010  (
            .Z (_N10183_2441),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I4)|(~I1&~I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7011  */ #(
            .INIT(32'b10111001000111010111100001000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7011  (
            .Z (_N10183_2442),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I4)|(~I0&I1&~I2&~I3)|(I0&I1&~I2&I3)|(~I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7024  */ #(
            .INIT(32'b11001100111111101010111010100011))
        \u_lcd_rgb_char/u_lcd_display/N9971_7024  (
            .Z (_N10183_2455),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&~I2&~I3&~I4)|(I0&~I1&~I4)|(I2&~I3&I4)|(I1&I4)|(I0&~I1&~I3)|(I1&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7025  */ #(
            .INIT(32'b11110010001100111111101111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7025  (
            .Z (_N10183_2456),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I3&~I4)|(~I1&I3&~I4)|(I0&~I4)|(~I1&~I3&I4)|(I2&I3)|(~I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7026  */ #(
            .INIT(32'b11111110111111101110111000010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7026  (
            .Z (_N10183_2457),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I2&I4)|(I0&I4)|(I1&I3)|(I0&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7027  */ #(
            .INIT(32'b10110011001101111111101100001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_7027  (
            .Z (_N10183_2458),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&~I2&~I4)|(~I0&~I2&~I3&I4)|(~I1&I4)|(I0&I2&I3)|(~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7028  */ #(
            .INIT(32'b11111011111111111111101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_7028  (
            .Z (_N10183_2459),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I3&I4)|(I2)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7029  */ #(
            .INIT(32'b10111011101110111111101110011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_7029  (
            .Z (_N10183_2460),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&I4)|(I0&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7053  */ #(
            .INIT(32'b10111111101111111101010101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7053  (
            .Z (_N10183_2484),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I4)|(I0&I4)|(~I2&~I3)|(I0&I1&I2&I3)|(~I0&~I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7055  */ #(
            .INIT(32'b10100101101001010100000001001111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7055  (
            .Z (_N10183_2486),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I4)|(I0&I2&I4) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_7060  */ #(
            .INIT(16'b1011111110110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7060  (
            .Z (_N10183_2491),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3)|(~I0&~I2)|(I0&I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7072  */ #(
            .INIT(32'b11101101111111011010110001010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7072  (
            .Z (_N10183_2503),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(I0&I2&I3)|(I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7075  */ #(
            .INIT(32'b11101101111111010101010111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7075  (
            .Z (_N10183_2506),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I3&~I4)|(~I0&~I4)|(I0&I2&I4)|(I1&I4)|(~I0&~I3)|(~I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7076  */ #(
            .INIT(32'b10101011111011111011100110111001))
        \u_lcd_rgb_char/u_lcd_display/N9971_7076  (
            .Z (_N10183_2507),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I4)|(I1&~I3&I4)|(I0&I4)|(~I0&~I1&~I2)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7077  */ #(
            .INIT(32'b10111010001000100100011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_7077  (
            .Z (_N10183_2508),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I2&~I3&~I4)|(~I0&I1&I3&~I4)|(~I1&I2&I3&I4)|(I0&I3&I4)|(I0&~I1&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7078  */ #(
            .INIT(32'b11111111111101111110111111011110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7078  (
            .Z (_N10183_2509),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(~I1&I4)|(~I0&I2&~I3)|(~I2&I3)|(I0&I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7080  */ #(
            .INIT(32'b11100101111111111011101011101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7080  (
            .Z (_N10183_2511),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I1&I2&I3&~I4)|(I0&~I4)|(~I3&I4)|(~I0&~I2&I4)|(~I0&I1&I4)|(I1&~I3)|(I0&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7081  */ #(
            .INIT(32'b10111001110111101111111111001110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7081  (
            .Z (_N10183_2512),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I2&~I4)|(I1&~I4)|(~I0&~I1&I2&I4)|(I0&~I2&~I3)|(I1&~I3)|(I0&I2&I3)|(~I0&~I1&I3)|(I0&I1) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_7082_3  */ #(
            .INIT(16'b1111111111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7082_3  (
            .Z (_N10183_2513),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7083  */ #(
            .INIT(32'b11111111111110111111101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7083  (
            .Z (_N10183_2514),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(~I1&I3)|(~I1&~I2)|(I1&I2)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7084  */ #(
            .INIT(32'b10011010100100111110101111101001))
        \u_lcd_rgb_char/u_lcd_display/N9971_7084  (
            .Z (_N10183_2515),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I2&~I4)|(I1&I2&~I4)|(I0&I2&~I4)|(I0&I1&~I4)|(I0&~I1&~I2&I4)|(~I0&~I1&I2&I4)|(~I0&~I1&~I2&~I3)|(I0&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7085  */ #(
            .INIT(32'b11111101111011110000011010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_7085  (
            .Z (_N10183_2516),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(I0&~I3&I4)|(~I0&I3&I4)|(~I0&~I2&I4)|(I0&I2&I4)|(I1&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7086  */ #(
            .INIT(32'b11110111111111010000010010000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_7086  (
            .Z (_N10183_2517),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&I4)|(~I1&I3&I4)|(I2&I4)|(~I0&I4)|(I0&I1&I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7089  */ #(
            .INIT(32'b11001001110001000000001100001101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7089  (
            .Z (_N10183_2520),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(~I0&~I1&~I2&~I4)|(I0&I1&I3&I4)|(I1&I2&I4)|(~I0&I1&~I2&~I3)|(~I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7108  */ #(
            .INIT(32'b11001100000000010001011000000001))
        \u_lcd_rgb_char/u_lcd_display/N9971_7108  (
            .Z (_N10183_2539),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I0&~I1&I2&I3&~I4)|(I1&I3&I4)|(~I0&~I1&~I2&~I3)|(~I0&I1&~I2&I3) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_7117  */ #(
            .INIT(4'b1001))
        \u_lcd_rgb_char/u_lcd_display/N9971_7117  (
            .Z (_N10183_2548),
            .I0 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = ~I1^I0 ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7138  */ #(
            .INIT(32'b11011111101010111111111010111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7138  (
            .Z (_N10183_2569),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I2&~I4)|(~I1&I2&~I4)|(~I1&~I2&I4)|(~I1&~I2&~I3)|(I0&~I3)|(~I0&I2&I3)|(I1&I3)|(I0&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7139  */ #(
            .INIT(32'b11111111010111101110010010101110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7139  (
            .Z (_N10183_2570),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I2&~I4)|(I3&I4)|(~I0&I2&I4)|(I0&~I2&~I3)|(~I0&I1&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7140  */ #(
            .INIT(32'b11110010000000001000101100010000))
        \u_lcd_rgb_char/u_lcd_display/N9971_7140  (
            .Z (_N10183_2571),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&I2&~I3&~I4)|(~I1&~I2&I3&~I4)|(I0&I1&I3&~I4)|(I2&I3&I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7141  */ #(
            .INIT(32'b10010000011001101001000101100100))
        \u_lcd_rgb_char/u_lcd_display/N9971_7141  (
            .Z (_N10183_2572),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&I3&~I4)|(I0&~I1&~I3&I4)|(I0&~I1&I2&~I3)|(~I0&I1&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7146  */ #(
            .INIT(32'b11111111110111111111101111011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7146  (
            .Z (_N10183_2577),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7147  */ #(
            .INIT(32'b11111110111111111101011011110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7147  (
            .Z (_N10183_2578),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&I4)|(~I1&~I3)|(I0&~I1&~I2)|(I1&I2)|(~I0&I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7148  */ #(
            .INIT(32'b10111001000111010111100001000110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7148  (
            .Z (_N10183_2579),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I1&~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(I0&I1&I3&I4)|(I0&I1&~I2&I4)|(~I0&~I1&I4)|(~I0&I1&~I2&~I3)|(I0&I1&~I2&I3)|(~I1&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7161  */ #(
            .INIT(32'b11001100111111101010111010100011))
        \u_lcd_rgb_char/u_lcd_display/N9971_7161  (
            .Z (_N10183_2592),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I1&~I2&~I3&~I4)|(I0&~I1&~I4)|(I2&~I3&I4)|(I1&I4)|(I0&~I1&~I3)|(I1&~I2&I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7162  */ #(
            .INIT(32'b11110010001100111111101111111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7162  (
            .Z (_N10183_2593),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I3&~I4)|(~I1&I3&~I4)|(I0&~I4)|(~I1&~I3&I4)|(I2&I3)|(~I1&I2)|(I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7163  */ #(
            .INIT(32'b11111110111111101110111000010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7163  (
            .Z (_N10183_2594),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I2&I4)|(I0&I4)|(I1&I3)|(I0&I3)|(~I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7164  */ #(
            .INIT(32'b10110011001101111111101100001010))
        \u_lcd_rgb_char/u_lcd_display/N9971_7164  (
            .Z (_N10183_2595),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&~I2&~I4)|(~I0&~I2&~I3&I4)|(~I1&I4)|(I0&I2&I3)|(~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7165  */ #(
            .INIT(32'b11111011111111111111101111111011))
        \u_lcd_rgb_char/u_lcd_display/N9971_7165  (
            .Z (_N10183_2596),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I3&I4)|(I2)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7166  */ #(
            .INIT(32'b10111011101110111111101110011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_7166  (
            .Z (_N10183_2597),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&I3&~I4)|(I0&I4)|(I0&I3)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7190  */ #(
            .INIT(32'b10111111101111111101010101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7190  (
            .Z (_N10183_2621),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I4)|(I0&I4)|(~I2&~I3)|(I0&I1&I2&I3)|(~I0&~I2)|(~I0&~I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_7192  */ #(
            .INIT(32'b10100101101001010100000001001111))
        \u_lcd_rgb_char/u_lcd_display/N9971_7192  (
            .Z (_N10183_2623),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&I1&I2&~I4)|(~I0&~I2&I4)|(I0&I2&I4) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_7197  */ #(
            .INIT(16'b1011111110110101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7197  (
            .Z (_N10183_2628),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3)|(~I0&~I2)|(I0&I2)|(~I0&~I1) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_7211  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7211  (
            .Z (_N10183_2642),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_7219  */ #(
            .INIT(4'b1101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7219  (
            .Z (_N10183_2650),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1)|(~I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_7279  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7279  (
            .Z (_N10183_2710),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_7281  */ #(
            .INIT(8'b11010100))
        \u_lcd_rgb_char/u_lcd_display/N9971_7281  (
            .Z (_N10183_2712),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&I2)|(~I0&I2)|(~I0&I1) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_7289  */ #(
            .INIT(4'b1001))
        \u_lcd_rgb_char/u_lcd_display/N9971_7289  (
            .Z (_N10183_2720),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ));
	// LUT = ~I1^I0 ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_7351  */ #(
            .INIT(16'b1011000100010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7351  (
            .Z (_N10183_2782),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&~I3)|(I0&I2&I3)|(~I0&~I1) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_7359  */ #(
            .INIT(8'b11000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_7359  (
            .Z (_N10183_2790),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I0&~I1&~I2)|(I1&I2) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_7421  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7421  (
            .Z (_N10183_2852),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_7480  */ #(
            .INIT(16'b1011000100010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7480  (
            .Z (_N10183_2911),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&~I3)|(I0&I2&I3)|(~I0&~I1) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_7545  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7545  (
            .Z (_N10183_2976),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_7601  */ #(
            .INIT(16'b1011000100010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7601  (
            .Z (_N10183_3032),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&~I3)|(I0&I2&I3)|(~I0&~I1) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_7666  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7666  (
            .Z (_N10183_3097),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_7722  */ #(
            .INIT(16'b1011000100010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7722  (
            .Z (_N10183_3153),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&~I3)|(I0&I2&I3)|(~I0&~I1) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_7787  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7787  (
            .Z (_N10183_3218),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_7843  */ #(
            .INIT(16'b1011000100010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7843  (
            .Z (_N10183_3274),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&~I3)|(I0&I2&I3)|(~I0&~I1) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_7908  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_7908  (
            .Z (_N10183_3339),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_7964  */ #(
            .INIT(16'b1011000100010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_7964  (
            .Z (_N10183_3395),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&~I3)|(I0&I2&I3)|(~I0&~I1) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_8029  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_8029  (
            .Z (_N10183_3460),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_display/N9971_8085  */ #(
            .INIT(16'b1011000100010101))
        \u_lcd_rgb_char/u_lcd_display/N9971_8085  (
            .Z (_N10183_3516),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I0&~I2&~I3)|(I0&I2&I3)|(~I0&~I1) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_8125  */ #(
            .INIT(4'b1011))
        \u_lcd_rgb_char/u_lcd_display/N9971_8125  (
            .Z (_N10183_3556),
            .I0 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I1)|(I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_8555  */ #(
            .INIT(8'b11111110))
        \u_lcd_rgb_char/u_lcd_display/N9971_8555  (
            .Z (_N10456),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_8566  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_8566  (
            .Z (_N10495),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_8567  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_8567  (
            .Z (_N10496),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_8570  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_8570  (
            .Z (_N10499),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_8571  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_8571  (
            .Z (_N10500),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_8572  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_8572  (
            .Z (_N10501),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_8573  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_8573  (
            .Z (_N10502),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_8575  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_8575  (
            .Z (_N10505),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1)|(I0) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_8681  (
            .Z (_N10183_1051),
            .I0 (_N10911_3),
            .I1 (_N10911_2),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_8780  */ #(
            .INIT(32'b10000011100000011110111111100011))
        \u_lcd_rgb_char/u_lcd_display/N9971_8780  (
            .Z (_N10924_2),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1&I3&~I4)|(I1&I2&~I4)|(I0&~I1&~I4)|(~I1&~I2&I3)|(~I0&~I1&~I2)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_8874  */ #(
            .INIT(32'b10111010110111111111111101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_8874  (
            .Z (_N10183_2373),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I4)|(I0&I1&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_8960  */ #(
            .INIT(32'b10111010110111111111111101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_8960  (
            .Z (_N10183_2099),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I4)|(I0&I1&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_9557  */ #(
            .INIT(32'b11100000000001001110000001011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_9557  (
            .Z (_N11004_2),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&~I3&~I4)|(~I0&I1&~I2&~I3)|(I1&I2&I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_9573  */ #(
            .INIT(32'b11110000000000011111111011101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_9573  (
            .Z (_N10183_1488),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(I0&~I4)|(~I0&~I1&~I2&~I3)|(I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_9710  */ #(
            .INIT(32'b11100000000001001110000001011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_9710  (
            .Z (_N11016_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&~I3&~I4)|(~I0&I1&~I2&~I3)|(I1&I2&I3)|(I0&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_9951  (
            .Z (_N10183_1326),
            .I0 (_N11036_3),
            .I1 (_N11036_2),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_9995  */ #(
            .INIT(32'b10111010110111111111111101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_9995  (
            .Z (_N10183_2236),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I4)|(I0&I1&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_10148  */ #(
            .INIT(32'b10111010110111111111111101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_10148  (
            .Z (_N10183_1962),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I4)|(I0&I1&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_10227  */ #(
            .INIT(32'b10111010110111111111111101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_10227  (
            .Z (_N10183_1825),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I4)|(I0&I1&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_11580  */ #(
            .INIT(32'b11110000000000011111111011101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_11580  (
            .Z (_N10183_1031),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(I0&~I4)|(~I0&~I1&~I2&~I3)|(I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_11607  (
            .Z (_N10183_1235),
            .I0 (_N11162_3),
            .I1 (_N11162_2),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_11613  */ #(
            .INIT(32'b11110000000000011111111011101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_11613  (
            .Z (_N10183_1579),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(I0&~I4)|(~I0&~I1&~I2&~I3)|(I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_11624  */ #(
            .INIT(32'b11110000000000011111111011101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_11624  (
            .Z (_N10183_1397),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(I0&~I4)|(~I0&~I1&~I2&~I3)|(I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_11632  */ #(
            .INIT(32'b11100000000001001110000001011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_11632  (
            .Z (_N11168_2),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&~I3&~I4)|(~I0&I1&~I2&~I3)|(I1&I2&I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_11703  */ #(
            .INIT(32'b11100000000001001110000001011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_11703  (
            .Z (_N11179_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&~I3&~I4)|(~I0&I1&~I2&~I3)|(I1&I2&I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_11848  */ #(
            .INIT(32'b11100000000001001110000001011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_11848  (
            .Z (_N11190_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&~I3&~I4)|(~I0&I1&~I2&~I3)|(I1&I2&I3)|(I0&I2&I3) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_12246  (
            .Z (_N10183_1508),
            .I0 (_N11227_3),
            .I1 (_N11227_2),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_12552  (
            .Z (_N10183_1417),
            .I0 (_N11259_3),
            .I1 (_N11259_2),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_13400  */ #(
            .INIT(32'b11110000000000011111111011101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_13400  (
            .Z (_N11319_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(I0&~I4)|(~I0&~I1&~I2&~I3)|(I2&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_14479  */ #(
            .INIT(32'b11000101110001011010101011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_14479  (
            .Z (_N11364_2),
            .I0 (_N10183_534),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [7] ),
            .ID (_N10183_292));
	// LUT = (~I3&~I4)|(ID&~I4)|(~I0&~I2&I4)|(I1&I2&I4) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_15686  (
            .Z (_N10183_1144),
            .I0 (_N11428_3),
            .I1 (_N11428_2),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_16034  (
            .Z (_N10183_1599),
            .I0 (_N11482_3),
            .I1 (_N11482_2),
            .S (\u_lcd_rgb_char/pixel_xpos_w [0] ));

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_16064  */ #(
            .INIT(32'b11100000000001001110000001011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_16064  (
            .Z (_N11489_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&~I3&~I4)|(~I0&I1&~I2&~I3)|(I1&I2&I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_16186  */ #(
            .INIT(32'b11100000000001001110000001011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_16186  (
            .Z (_N11502_2),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (~I2&~I3&~I4)|(~I0&~I3&~I4)|(~I0&I1&~I2&~I3)|(I1&I2&I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_16192  */ #(
            .INIT(32'b11110000000000011111111011101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_16192  (
            .Z (_N11503_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(I0&~I4)|(~I0&~I1&~I2&~I3)|(I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_17128  */ #(
            .INIT(32'b11110000000000011111111011101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_17128  (
            .Z (_N10183_1215),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I1&~I4)|(I0&~I4)|(~I0&~I1&~I2&~I3)|(I2&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_17586  */ #(
            .INIT(32'b10111010110111111111111101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_17586  (
            .Z (_N10183_1675),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I4)|(I0&I1&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&~I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_19961  */ #(
            .INIT(32'b10111010110111111111111101011111))
        \u_lcd_rgb_char/u_lcd_display/N9971_19961  (
            .Z (_N10183_2510),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I4)|(I0&I1&I4)|(~I0&~I3)|(I0&I3)|(I0&~I2)|(~I0&~I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_display/N9971_20029  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_display/N9971_20029  (
            .Z (_N12065),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20033  */ #(
            .INIT(32'b11111111111111111111101111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20033  (
            .Z (_N10911_2),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I4)|(~I0&~I3)|(I0&I3)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20038  */ #(
            .INIT(32'b11111111111111111111101111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20038  (
            .Z (_N11428_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I4)|(~I0&~I3)|(I0&I3)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20043  */ #(
            .INIT(32'b11111111111111111111101111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20043  (
            .Z (_N11162_2),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I4)|(~I0&~I3)|(I0&I3)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20048  */ #(
            .INIT(32'b11111111111111111111101111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20048  (
            .Z (_N11036_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I4)|(~I0&~I3)|(I0&I3)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20053  */ #(
            .INIT(32'b11111111111111111111101111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20053  (
            .Z (_N11259_2),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I4)|(~I0&~I3)|(I0&I3)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20058  */ #(
            .INIT(32'b11111111111111111111101111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20058  (
            .Z (_N11227_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I4)|(~I0&~I3)|(I0&I3)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20063  */ #(
            .INIT(32'b11111111111111111111101111011101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20063  (
            .Z (_N11482_2),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I4)|(~I0&~I3)|(I0&I3)|(~I0&I2)|(~I0&~I1)|(I0&I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20157  */ #(
            .INIT(32'b10111111101011111111111101110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20157  (
            .Z (_N12282),
            .I0 (_N10495),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_2790),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I3&~I4)|(~I1&~I4)|(~ID&~I4)|(~I2&I4)|(I0&I4)|(~I1&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20159  */ #(
            .INIT(32'b10111111101011111111111101110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20159  (
            .Z (_N12284),
            .I0 (_N10496),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_2790),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I3&~I4)|(~I1&~I4)|(~ID&~I4)|(~I2&I4)|(I0&I4)|(~I1&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20161  */ #(
            .INIT(32'b10111111101011111111111101110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20161  (
            .Z (_N12286),
            .I0 (_N10502),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_2790),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I3&~I4)|(~I1&~I4)|(~ID&~I4)|(~I2&I4)|(I0&I4)|(~I1&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20163  */ #(
            .INIT(32'b10111111101011111111111101110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20163  (
            .Z (_N12288),
            .I0 (_N10499),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_2790),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I3&~I4)|(~I1&~I4)|(~ID&~I4)|(~I2&I4)|(I0&I4)|(~I1&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20165  */ #(
            .INIT(32'b10111111101011111111111101110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20165  (
            .Z (_N12290),
            .I0 (_N10505),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_2790),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I3&~I4)|(~I1&~I4)|(~ID&~I4)|(~I2&I4)|(I0&I4)|(~I1&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20167  */ #(
            .INIT(32'b10111111101011111111111101110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20167  (
            .Z (_N12292),
            .I0 (_N10500),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_2790),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I3&~I4)|(~I1&~I4)|(~ID&~I4)|(~I2&I4)|(I0&I4)|(~I1&I3) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20169  */ #(
            .INIT(32'b10111111101011111111111101110111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20169  (
            .Z (_N12294),
            .I0 (_N10501),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I2 (_N10183_2790),
            .I3 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (I3&~I4)|(~I1&~I4)|(~ID&~I4)|(~I2&I4)|(I0&I4)|(~I1&I3) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20171  */ #(
            .INIT(32'b11110101111101011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20171  (
            .Z (_N10183_1795),
            .I0 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I4)|(~I0&I4)|(~I0&~I3)|(I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20173  */ #(
            .INIT(32'b11110101111101011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20173  (
            .Z (_N10183_1935),
            .I0 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I4)|(~I0&I4)|(~I0&~I3)|(I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20175  */ #(
            .INIT(32'b11110101111101011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20175  (
            .Z (_N10183_2072),
            .I0 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I4)|(~I0&I4)|(~I0&~I3)|(I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20177  */ #(
            .INIT(32'b11110101111101011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20177  (
            .Z (_N10183_2209),
            .I0 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I4)|(~I0&I4)|(~I0&~I3)|(I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20179  */ #(
            .INIT(32'b11110101111101011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20179  (
            .Z (_N10183_2346),
            .I0 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I4)|(~I0&I4)|(~I0&~I3)|(I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20181  */ #(
            .INIT(32'b11110101111101011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20181  (
            .Z (_N10183_2483),
            .I0 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I4)|(~I0&I4)|(~I0&~I3)|(I2)|(~I0&I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20183  */ #(
            .INIT(32'b11110101111101011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20183  (
            .Z (_N10183_2620),
            .I0 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I0&~I4)|(~I0&I4)|(~I0&~I3)|(I2)|(~I0&I1) ;

    GTP_MUX2LUT6 \u_lcd_rgb_char/u_lcd_display/N9971_20199  (
            .Z (_N12317),
            .I0 (_N10183_174),
            .I1 (_N10183_306),
            .S (\u_lcd_rgb_char/pixel_xpos_w [1] ));

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_20217  */ #(
            .INIT(8'b11111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20217  (
            .Z (_N10183_2789),
            .I0 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(~I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_20221  */ #(
            .INIT(8'b11111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20221  (
            .Z (_N10183_2918),
            .I0 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(~I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_20225  */ #(
            .INIT(8'b11111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20225  (
            .Z (_N10183_3039),
            .I0 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(~I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_20229  */ #(
            .INIT(8'b11111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20229  (
            .Z (_N10183_3160),
            .I0 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(~I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_20233  */ #(
            .INIT(8'b11111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20233  (
            .Z (_N10183_3281),
            .I0 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(~I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_20237  */ #(
            .INIT(8'b11111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20237  (
            .Z (_N10183_3402),
            .I0 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(~I0) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_display/N9971_20241  */ #(
            .INIT(8'b11111101))
        \u_lcd_rgb_char/u_lcd_display/N9971_20241  (
            .Z (_N10183_3523),
            .I0 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I1 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I2)|(I1)|(~I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20320  */ #(
            .INIT(32'b11101011110000101100101111000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_20320  (
            .Z (_N10183_1686),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I1&~I2&I3)|(I0&I1&I3)|(I0&~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20335  */ #(
            .INIT(32'b11101011110000101100101111000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_20335  (
            .Z (_N10183_2247),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I1&~I2&I3)|(I0&I1&I3)|(I0&~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20340  */ #(
            .INIT(32'b11111111111110111111101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20340  (
            .Z (_N10183_2240),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(~I1&I3)|(~I1&~I2)|(I1&I2)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20365  */ #(
            .INIT(32'b11101011110000101100101111000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_20365  (
            .Z (_N10183_1973),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I1&~I2&I3)|(I0&I1&I3)|(I0&~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20370  */ #(
            .INIT(32'b11111111111110111111101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20370  (
            .Z (_N10183_1966),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(~I1&I3)|(~I1&~I2)|(I1&I2)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20375  */ #(
            .INIT(32'b11101011110000101100101111000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_20375  (
            .Z (_N10183_1836),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I1&~I2&I3)|(I0&I1&I3)|(I0&~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20380  */ #(
            .INIT(32'b11111111111110111111101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20380  (
            .Z (_N10183_1829),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(~I1&I3)|(~I1&~I2)|(I1&I2)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20415  */ #(
            .INIT(32'b11101011110000101100101111000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_20415  (
            .Z (_N10183_2384),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I1&~I2&I3)|(I0&I1&I3)|(I0&~I1&~I2)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20423  */ #(
            .INIT(32'b11111111111111011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20423  (
            .Z (_N10183_786),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [10] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (~I3&~I4)|(I3&I4)|(~I0&~I3)|(ID&I3)|(I2)|(I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20478  */ #(
            .INIT(32'b11111111111110111111101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20478  (
            .Z (_N10183_2377),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(~I1&I3)|(~I1&~I2)|(I1&I2)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20506  */ #(
            .INIT(32'b11101011110000101100101111000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_20506  (
            .Z (_N10183_2110),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I1&~I2&I3)|(I0&I1&I3)|(I0&~I1&~I2)|(I1&I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20511  */ #(
            .INIT(32'b11111111111110111111101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20511  (
            .Z (_N10183_2103),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(~I1&I3)|(~I1&~I2)|(I1&I2)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20619  */ #(
            .INIT(32'b10001010101010110000000000000000))
        \u_lcd_rgb_char/u_lcd_display/N9971_20619  (
            .Z (_N10183_956),
            .I0 (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .I1 (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_display/N59 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [6] ));
	// LUT = (~I1&~I2&~I3&I4)|(I0&~I3&I4)|(I0&~I2&I4)|(I0&I1&I4) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20661  */ #(
            .INIT(32'b11101110000010011110111011011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_20661  (
            .Z (_N10183_1743),
            .I0 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I1&I2&~I4)|(~I0&~I1&~I2&~I3)|(I1&I3)|(I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20736  */ #(
            .INIT(32'b11111111111110111111101111101111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20736  (
            .Z (_N10183_1679),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I1&~I3&~I4)|(I3&I4)|(~I1&I4)|(~I1&I3)|(~I1&~I2)|(I1&I2)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20770  */ #(
            .INIT(32'b11101110000010011110111011011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_20770  (
            .Z (_N10183_2299),
            .I0 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I1&I2&~I4)|(~I0&~I1&~I2&~I3)|(I1&I3)|(I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20818  */ #(
            .INIT(32'b11101110000010011110111011011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_20818  (
            .Z (_N10183_2573),
            .I0 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I1&I2&~I4)|(~I0&~I1&~I2&~I3)|(I1&I3)|(I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20823  */ #(
            .INIT(32'b11101110000010011110111011011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_20823  (
            .Z (_N10183_2162),
            .I0 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I1&I2&~I4)|(~I0&~I1&~I2&~I3)|(I1&I3)|(I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20845  */ #(
            .INIT(32'b11101110000010011110111011011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_20845  (
            .Z (_N10183_2025),
            .I0 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I1&I2&~I4)|(~I0&~I1&~I2&~I3)|(I1&I3)|(I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20880  */ #(
            .INIT(32'b11101110000010011110111011011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_20880  (
            .Z (_N10183_1888),
            .I0 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I1&I2&~I4)|(~I0&~I1&~I2&~I3)|(I1&I3)|(I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20909  */ #(
            .INIT(32'b11101110000010011110111011011001))
        \u_lcd_rgb_char/u_lcd_display/N9971_20909  (
            .Z (_N10183_2436),
            .I0 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (~I0&~I1&~I3&~I4)|(I1&I2&~I4)|(~I0&~I1&~I2&~I3)|(I1&I3)|(I0&I3)|(I0&I1&~I2) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20937  */ #(
            .INIT(32'b11101011110000101100101111000010))
        \u_lcd_rgb_char/u_lcd_display/N9971_20937  (
            .Z (_N10183_2521),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ));
	// LUT = (I0&I3&I4)|(~I1&~I2&I3)|(I0&I1&I3)|(I0&~I1&~I2)|(I1&I2) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20942  */ #(
            .INIT(32'b11111111111111011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20942  (
            .Z (_N10183_560),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (~I3&~I4)|(I3&I4)|(~I0&~I3)|(ID&I3)|(I2)|(I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20949  */ #(
            .INIT(32'b11111111111111011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20949  (
            .Z (_N10183_618),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [2] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (~I3&~I4)|(I3&I4)|(~I0&~I3)|(ID&I3)|(I2)|(I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20956  */ #(
            .INIT(32'b11111111111111011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20956  (
            .Z (_N10183_730),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [6] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (~I3&~I4)|(I3&I4)|(~I0&~I3)|(ID&I3)|(I2)|(I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20963  */ #(
            .INIT(32'b11111111111111011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20963  (
            .Z (_N10183_842),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [10] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (~I3&~I4)|(I3&I4)|(~I0&~I3)|(ID&I3)|(I2)|(I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20970  */ #(
            .INIT(32'b11111111111111011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20970  (
            .Z (_N10183_898),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I3 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I4 (\u_lcd_rgb_char/bcd_data_x [14] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (~I3&~I4)|(I3&I4)|(~I0&~I3)|(ID&I3)|(I2)|(I1) ;

    GTP_LUT5M /* \u_lcd_rgb_char/u_lcd_display/N9971_20977  */ #(
            .INIT(32'b11111111111111011111111011111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20977  (
            .Z (_N10183_674),
            .I0 (_N10183_1004),
            .I1 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I3 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I4 (\u_lcd_rgb_char/bcd_data_y [6] ),
            .ID (\u_lcd_rgb_char/pixel_xpos_w [0] ));
	// LUT = (~I3&~I4)|(I3&I4)|(~I0&~I3)|(ID&I3)|(I2)|(I1) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20990  */ #(
            .INIT(32'b10111011111111111111101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20990  (
            .Z (_N10911_3),
            .I0 (\u_lcd_rgb_char/bcd_data_y [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&~I4)|(~I3)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20993  */ #(
            .INIT(32'b10111011111111111111101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20993  (
            .Z (_N11428_3),
            .I0 (\u_lcd_rgb_char/bcd_data_x [0] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [1] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&~I4)|(~I3)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20996  */ #(
            .INIT(32'b10111011111111111111101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20996  (
            .Z (_N11162_3),
            .I0 (\u_lcd_rgb_char/bcd_data_y [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&~I4)|(~I3)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_20999  */ #(
            .INIT(32'b10111011111111111111101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_20999  (
            .Z (_N11036_3),
            .I0 (\u_lcd_rgb_char/bcd_data_x [4] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [5] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&~I4)|(~I3)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_21002  */ #(
            .INIT(32'b10111011111111111111101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_21002  (
            .Z (_N11259_3),
            .I0 (\u_lcd_rgb_char/bcd_data_y [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_y [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_y [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&~I4)|(~I3)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_21005  */ #(
            .INIT(32'b10111011111111111111101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_21005  (
            .Z (_N11227_3),
            .I0 (\u_lcd_rgb_char/bcd_data_x [8] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [9] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [11] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&~I4)|(~I3)|(~I1)|(I0) ;

    GTP_LUT5 /* \u_lcd_rgb_char/u_lcd_display/N9971_21008  */ #(
            .INIT(32'b10111011111111111111101111111111))
        \u_lcd_rgb_char/u_lcd_display/N9971_21008  (
            .Z (_N11482_3),
            .I0 (\u_lcd_rgb_char/bcd_data_x [12] ),
            .I1 (\u_lcd_rgb_char/bcd_data_x [13] ),
            .I2 (\u_lcd_rgb_char/bcd_data_x [15] ),
            .I3 (\u_lcd_rgb_char/u_lcd_display/N59 [5] ),
            .I4 (\u_lcd_rgb_char/u_lcd_display/N59 [8] ));
	// LUT = (I2&~I4)|(~I3)|(~I1)|(I0) ;

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_display/pixel_data[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_display/pixel_data[0]  (
            .Q (\u_lcd_rgb_char/pixel_data_w [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_display/N9971 [0] ));
	// ../../rtl/lcd_rgb_char/lcd_display.v:117

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N0  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_driver/N0  (
            .Z (\u_lcd_rgb_char/lcd_rgb_o [0] ),
            .I0 (nt_lcd_de),
            .I1 (\u_lcd_rgb_char/pixel_data_w [0] ));
	// LUT = I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:127

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_0  */ #(
            .INIT(32'b11111111111111110000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [0] ),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b1 ;
	// CARRY = (1'b0) ? CIN : (1'b1) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_1  */ #(
            .INIT(32'b01101001011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [1] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [0] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [0] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [0] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [0] ),
            .ID ());
	// LUT = ~I2^I1^CIN ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_2  */ #(
            .INIT(32'b01101001011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [2] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [1] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [1] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_cnt[1]_inv ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_cnt[1]_inv ),
            .ID ());
	// LUT = ~I2^I1^CIN ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_3  */ #(
            .INIT(32'b01101001011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [3] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [2] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [2] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb0 [2] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb0 [2] ),
            .ID ());
	// LUT = ~I2^I1^CIN ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_4  */ #(
            .INIT(32'b01011010011010011111000011000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [4] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [3] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [3] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb0 [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb0 [3] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(CIN&~I2&I3)|(~CIN&I2&I3)|(CIN&I1&~I2)|(~CIN&I1&I2) ;
	// CARRY = ((~I1&~I2&~I3)|(I2&I3)|(I1&I2)) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_5  */ #(
            .INIT(32'b01101001011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_5  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [5] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [4] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [4] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb0 [4] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb0 [4] ),
            .ID ());
	// LUT = ~I2^I1^CIN ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_6  */ #(
            .INIT(32'b01101001011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_6  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [6] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [5] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [5] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb0 [5] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb0 [5] ),
            .ID ());
	// LUT = ~I2^I1^CIN ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_7  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_7  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [7] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [6] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [6] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb0 [6] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb0 [6] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_8  */ #(
            .INIT(32'b01101001011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_8  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [8] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [7] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [7] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb0 [7] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb0 [7] ),
            .ID ());
	// LUT = ~I2^I1^CIN ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_9  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_9  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [9] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [8] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [8] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb0 [8] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb0 [8] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_10  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_10  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [10] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [9] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [9] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb0 [9] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb0 [9] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_11  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_1.fsub_11  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb1 [10] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_1.co [10] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb0 [10] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb0 [10] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_0  */ #(
            .INIT(32'b11001100110011000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_0  (
            .COUT (_N690),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [1] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I1 ;
	// CARRY = (1'b0) ? CIN : (I1) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_1  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_1  (
            .COUT (_N691),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb0 [2] ),
            .CIN (_N690),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [2] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_2  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_2  (
            .COUT (_N692),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb0 [3] ),
            .CIN (_N691),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [3] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_3  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_3  (
            .COUT (_N693),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb0 [4] ),
            .CIN (_N692),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [4] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_4  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_4  (
            .COUT (_N694),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb0 [5] ),
            .CIN (_N693),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [5] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_5  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_5  (
            .COUT (_N695),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb0 [6] ),
            .CIN (_N694),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [6] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_6  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_6  (
            .COUT (_N696),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb0 [7] ),
            .CIN (_N695),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [7] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_7  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_7  (
            .COUT (_N697),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb0 [8] ),
            .CIN (_N696),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [8] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_8  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_8  (
            .COUT (_N698),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb0 [9] ),
            .CIN (_N697),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [9] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_3_9  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_3_9  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb0 [10] ),
            .CIN (_N698),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [10] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_0  */ #(
            .INIT(32'b11111111111111110000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [0] ),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b1 ;
	// CARRY = (1'b0) ? CIN : (1'b1) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_1  */ #(
            .INIT(32'b01101001000000001100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [1] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [1] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [0] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb1 [1] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [1] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&I3)|(CIN&I1&~I2&I3)|(CIN&~I1&I2&I3)|(~CIN&I1&I2&I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_2  */ #(
            .INIT(32'b01101001000000001100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [2] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [2] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [1] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb1 [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [2] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&I3)|(CIN&I1&~I2&I3)|(CIN&~I1&I2&I3)|(~CIN&I1&I2&I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_3  */ #(
            .INIT(32'b10010110000000000011110000111100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [3] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [3] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [2] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb1 [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [3] ),
            .ID ());
	// LUT = (CIN&~I1&~I2&I3)|(~CIN&I1&~I2&I3)|(~CIN&~I1&I2&I3)|(CIN&I1&I2&I3) ;
	// CARRY = (I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_4  */ #(
            .INIT(32'b01101001000000001100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [4] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [4] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [3] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb1 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [4] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&I3)|(CIN&I1&~I2&I3)|(CIN&~I1&I2&I3)|(~CIN&I1&I2&I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_5  */ #(
            .INIT(32'b10010000100100000011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_5  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [5] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [5] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [4] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb1 [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [5] ),
            .ID ());
	// LUT = (~CIN&~I1&I2)|(CIN&I1&I2) ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_6  */ #(
            .INIT(32'b01101001000000001100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_6  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [6] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [6] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [5] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb1 [6] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [6] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&I3)|(CIN&I1&~I2&I3)|(CIN&~I1&I2&I3)|(~CIN&I1&I2&I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_7  */ #(
            .INIT(32'b01101001000000001100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_7  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [7] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [7] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [6] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/nb1 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [7] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&I3)|(CIN&I1&~I2&I3)|(CIN&~I1&I2&I3)|(~CIN&I1&I2&I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_8  */ #(
            .INIT(32'b10010000100100000011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_8  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [8] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [8] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [7] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb1 [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [8] ),
            .ID ());
	// LUT = (~CIN&~I1&I2)|(CIN&I1&I2) ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_9  */ #(
            .INIT(32'b10010000100100000011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_9  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [9] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [9] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [8] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb1 [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [9] ),
            .ID ());
	// LUT = (~CIN&~I1&I2)|(CIN&I1&I2) ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_10  */ #(
            .INIT(32'b10010000100100000011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N7_4.fsub_10  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [10] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N7_4.co [9] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb1 [10] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb1 [10] ),
            .ID ());
	// LUT = (~CIN&~I1&I2)|(CIN&I1&I2) ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N12_1_0  */ #(
            .INIT(32'b00000000000000000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N12_1_0  (
            .COUT (_N619),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = (1'b0) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N12_1_1  */ #(
            .INIT(32'b10010110100101100011110000111100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N12_1_1  (
            .COUT (_N620),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N12 [0] ),
            .CIN (_N619),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [10] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .ID ());
	// LUT = I2^I1^CIN ;
	// CARRY = (I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N12_1_2  */ #(
            .INIT(32'b10101001101010010000001100000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N12_1_2  (
            .COUT (_N621),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N12 [1] ),
            .CIN (_N620),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I3 (),
            .I4 (1'b1),
            .ID ());
	// LUT = (~CIN&~I1&~I2)|(CIN&I2)|(CIN&I1) ;
	// CARRY = (~I1&~I2) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N12_1_3  */ #(
            .INIT(32'b01100110011001011100110011001111), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N12_1_3  (
            .COUT (_N622),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N12 [2] ),
            .CIN (_N621),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_clk_div/N39 ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .I4 (1'b0),
            .ID ());
	// LUT = (~CIN&~I2&~I3)|(CIN&~I1&I3)|(CIN&~I1&I2)|(~CIN&I1) ;
	// CARRY = ((~I2&~I3)|(I1)) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N12_1_4  */ #(
            .INIT(32'b10010110100101100011110000111100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N12_1_4  (
            .COUT (_N623),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N12 [3] ),
            .CIN (_N622),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .ID ());
	// LUT = I2^I1^CIN ;
	// CARRY = (I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N12_1_5  */ #(
            .INIT(32'b01100110011001011100110011001111), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N12_1_5  (
            .COUT (_N624),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N12 [4] ),
            .CIN (_N623),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_clk_div/N39 ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .I4 (1'b0),
            .ID ());
	// LUT = (~CIN&~I2&~I3)|(CIN&~I1&I3)|(CIN&~I1&I2)|(~CIN&I1) ;
	// CARRY = ((~I2&~I3)|(I1)) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N12_1_6  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N12_1_6  (
            .COUT (_N625),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N12 [5] ),
            .CIN (_N624),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N12_1_7  */ #(
            .INIT(32'b10101010101010100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N12_1_7  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N12 [6] ),
            .CIN (_N625),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = CIN ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N13.lt_0  */ #(
            .INIT(32'b00100000111100100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N13.lt_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N13.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N12 [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N12 [1] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [1] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = (1'b0) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N13.lt_1  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N13.lt_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N13.co [2] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N13.co [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N12 [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N12 [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [3] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N13.lt_2  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N13.lt_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N13.co [4] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N13.co [2] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N12 [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N12 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [5] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N13.lt_3  */ #(
            .INIT(32'b00000010000000100000100100001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N13.lt_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N13.co [6] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N13.co [4] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N12 [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [7] ),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I0&~I1&~I2 ;
	// CARRY = ((~I0&~I1&~I2)|(I0&I1&~I2)) ? CIN : (I0&~I1&~I2) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N13.lt_4  */ #(
            .INIT(32'b00000000000000000001000100010001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N13.lt_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N13.co [8] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N13.co [6] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [9] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = (~I0&~I1) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N13.lt_5  */ #(
            .INIT(32'b00100010001000100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N13.lt_5  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N13.co [8] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [10] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = CIN&~I1 ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N16_1_0  */ #(
            .INIT(32'b00000000000000000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N16_1_0  (
            .COUT (_N627),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = (1'b0) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N16_1_1  */ #(
            .INIT(32'b10010110100101100011110000111100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N16_1_1  (
            .COUT (_N628),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N16 [3] ),
            .CIN (_N627),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N12 [3] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N12 [3] ),
            .ID ());
	// LUT = I2^I1^CIN ;
	// CARRY = (I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N16_1_2  */ #(
            .INIT(32'b10100101100101100000111100111100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N16_1_2  (
            .COUT (_N629),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N16 [4] ),
            .CIN (_N628),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N12 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N12 [4] ),
            .ID ());
	// LUT = (CIN&~I1&~I2&~I3)|(~CIN&~I1&I2&~I3)|(~CIN&~I2&I3)|(CIN&I2&I3)|(~CIN&I1&~I2)|(CIN&I1&I2) ;
	// CARRY = ((~I1&I2&~I3)|(~I2&I3)|(I1&~I2)) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N16_1_3  */ #(
            .INIT(32'b10100101100101100000111100111100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N16_1_3  (
            .COUT (_N630),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N16 [5] ),
            .CIN (_N629),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N12 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N12 [5] ),
            .ID ());
	// LUT = (CIN&~I1&~I2&~I3)|(~CIN&~I1&I2&~I3)|(~CIN&~I2&I3)|(CIN&I2&I3)|(~CIN&I1&~I2)|(CIN&I1&I2) ;
	// CARRY = ((~I1&I2&~I3)|(~I2&I3)|(I1&~I2)) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N16_1_4  */ #(
            .INIT(32'b01011010011010011111000011000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N16_1_4  (
            .COUT (_N631),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N16 [6] ),
            .CIN (_N630),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N12 [6] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N12 [6] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(CIN&~I2&I3)|(~CIN&I2&I3)|(CIN&I1&~I2)|(~CIN&I1&I2) ;
	// CARRY = ((~I1&~I2&~I3)|(I2&I3)|(I1&I2)) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N16_1_5  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N16_1_5  (
            .COUT (_N632),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N16 [7] ),
            .CIN (_N631),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N16_1_6  */ #(
            .INIT(32'b10011001100110100011001100110000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N16_1_6  (
            .COUT (_N633),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N16 [8] ),
            .CIN (_N632),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_clk_div/N39 ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I2&~I3)|(~CIN&~I1&I3)|(~CIN&~I1&I2)|(CIN&I1) ;
	// CARRY = ((~I1&I3)|(~I1&I2)) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N16_1_7  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N16_1_7  (
            .COUT (_N634),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N16 [9] ),
            .CIN (_N633),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [10] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N16_1_8  */ #(
            .INIT(32'b10101010101010100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N16_1_8  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N16 [10] ),
            .CIN (_N634),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = CIN ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N17.lt_0  */ #(
            .INIT(32'b00100000111100100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N17.lt_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N17.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N12 [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N12 [1] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [1] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = (1'b0) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N17.lt_1  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N17.lt_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N17.co [2] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N17.co [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N12 [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N16 [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [3] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N17.lt_2  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N17.lt_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N17.co [4] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N17.co [2] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N16 [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N16 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [5] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N17.lt_3  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N17.lt_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N17.co [6] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N17.co [4] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N16 [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N16 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [7] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N17.lt_4  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N17.lt_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N17.co [8] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N17.co [6] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N16 [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N16 [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [9] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N17.lt_5  */ #(
            .INIT(32'b10100000111110100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N17.lt_5  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N17.co [8] ),
            .I0 (),
            .I1 (),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N16 [10] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [10] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(CIN&~I3)|(CIN&I2) ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:143

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_0  */ #(
            .INIT(32'b11001100110011000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_0  (
            .COUT (_N700),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [0] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I1 ;
	// CARRY = (1'b0) ? CIN : (I1) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_1  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_1  (
            .COUT (_N701),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [1] ),
            .CIN (_N700),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [1] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_2  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_2  (
            .COUT (_N702),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [2] ),
            .CIN (_N701),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [2] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_3  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_3  (
            .COUT (_N703),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [3] ),
            .CIN (_N702),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [3] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_4  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_4  (
            .COUT (_N704),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [4] ),
            .CIN (_N703),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [4] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_5  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_5  (
            .COUT (_N705),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [5] ),
            .CIN (_N704),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [5] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_6  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_6  (
            .COUT (_N706),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [6] ),
            .CIN (_N705),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [6] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_7  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_7  (
            .COUT (_N707),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [7] ),
            .CIN (_N706),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [7] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_8  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_8  (
            .COUT (_N708),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [8] ),
            .CIN (_N707),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [8] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_9  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_9  (
            .COUT (_N709),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [9] ),
            .CIN (_N708),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [9] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N23_1_10  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N23_1_10  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N23 [10] ),
            .CIN (_N709),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [10] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_0  */ #(
            .INIT(32'b11111111111111110000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [0] ),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b1 ;
	// CARRY = (1'b0) ? CIN : (1'b1) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_1  */ #(
            .INIT(32'b00000000011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [1] ),
            .Z (_N12225),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [0] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N12 [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/v_cnt[0]_inv ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/v_cnt[0]_inv ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(~CIN&I1&I2&~I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_2  */ #(
            .INIT(32'b00000000011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [2] ),
            .Z (_N12226),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [1] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N12 [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N23 [1] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [1] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(~CIN&I1&I2&~I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_3  */ #(
            .INIT(32'b00000000011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [3] ),
            .Z (_N12227),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [2] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N12 [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N23 [2] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [2] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(~CIN&I1&I2&~I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_4  */ #(
            .INIT(32'b00000000011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [4] ),
            .Z (_N12228),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [3] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N12 [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N23 [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [3] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(~CIN&I1&I2&~I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_5  */ #(
            .INIT(32'b00000000011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_5  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [5] ),
            .Z (_N12229),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [4] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N12 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N23 [4] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [4] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(~CIN&I1&I2&~I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_6  */ #(
            .INIT(32'b00000000011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_6  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [6] ),
            .Z (_N12230),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [5] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N12 [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N23 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [5] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(~CIN&I1&I2&~I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_7  */ #(
            .INIT(32'b00000000011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_7  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [7] ),
            .Z (_N12231),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [6] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N12 [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N23 [6] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [6] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(~CIN&I1&I2&~I3) ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_8  */ #(
            .INIT(32'b00001001000000000011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_8  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [8] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [7] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [7] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [7] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [7] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&I3)|(CIN&I1&~I2&I3) ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_9  */ #(
            .INIT(32'b00001001000000000011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_9  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [9] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [8] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [8] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [8] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&I3)|(CIN&I1&~I2&I3) ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_10  */ #(
            .INIT(32'b00001001000000000011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_10  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N25.co [10] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [9] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [9] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [9] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&I3)|(CIN&I1&~I2&I3) ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N25.fsub_11  */ #(
            .INIT(32'b00001001000000000011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N25.fsub_11  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [10] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N25.co [10] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [10] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N23 [10] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&I3)|(CIN&I1&~I2&I3) ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:144

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N98_1_0  */ #(
            .INIT(32'b00000000000000000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N98_1_0  (
            .COUT (_N636),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = (1'b0) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N98_1_1  */ #(
            .INIT(32'b10010110100101100011110000111100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N98_1_1  (
            .COUT (_N637),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N98 [1] ),
            .CIN (_N636),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .ID ());
	// LUT = I2^I1^CIN ;
	// CARRY = (I2^I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N98_1_2  */ #(
            .INIT(32'b10101010101010100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N98_1_2  (
            .COUT (_N638),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N98 [2] ),
            .CIN (_N637),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .ID ());
	// LUT = CIN ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N98_1_3  */ #(
            .INIT(32'b01010101010101011111111111111111), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N98_1_3  (
            .COUT (_N639),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N98 [3] ),
            .CIN (_N638),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = ~CIN ;
	// CARRY = (1'b1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N98_1_4  */ #(
            .INIT(32'b10011001100101100011001100111100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N98_1_4  (
            .COUT (_N640),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N98 [4] ),
            .CIN (_N639),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .ID ());
	// LUT = (CIN&~I1&~I2&~I3)|(~CIN&I1&~I2&~I3)|(~CIN&~I1&I3)|(CIN&I1&I3)|(~CIN&~I1&I2)|(CIN&I1&I2) ;
	// CARRY = ((I1&~I2&~I3)|(~I1&I3)|(~I1&I2)) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N98_1_5  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N98_1_5  (
            .COUT (_N641),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N98 [5] ),
            .CIN (_N640),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N98_1_6  */ #(
            .INIT(32'b01010110010101101111110011111100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N98_1_6  (
            .COUT (_N642),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N98 [6] ),
            .CIN (_N641),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I2)|(~CIN&I1) ;
	// CARRY = ((I2)|(I1)) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N98_1_7  */ #(
            .INIT(32'b10010110100101010011110000111111), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N98_1_7  (
            .COUT (_N643),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N98 [7] ),
            .CIN (_N642),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (\u_lcd_rgb_char/u_clk_div/N39 ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .ID ());
	// LUT = (~CIN&~I1&~I3)|(CIN&~I1&~I2&I3)|(~CIN&I1&~I2)|(~CIN&~I1&I2)|(CIN&I1&I2) ;
	// CARRY = ((~I1&~I3)|(I1&~I2)|(~I1&I2)) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N98_1_8  */ #(
            .INIT(32'b10101010101010100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N98_1_8  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N98 [8] ),
            .CIN (_N643),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = CIN ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_0  */ #(
            .INIT(32'b10101010101010100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N98 [1] ),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I0 ;
	// CARRY = (1'b0) ? CIN : (I0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_1  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [1] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N100 [2] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [0] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [2] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [2] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_2  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [2] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N100 [3] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [1] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [3] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [3] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_3  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [3] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N100 [4] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [2] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [4] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [4] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_4  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [4] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N100 [5] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [3] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [5] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [5] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_5  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_5  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [5] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N100 [6] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [4] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [6] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [6] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_6  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_6  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [6] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N100 [7] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [5] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [7] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [7] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_7  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_7  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [7] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N100 [8] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [6] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [8] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [8] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_8  */ #(
            .INIT(32'b01010101010101011111111111111111), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N100_1.fsub_8  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N100 [9] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N100_1.co [7] ),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~CIN ;
	// CARRY = (1'b1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N101.lt_0  */ #(
            .INIT(32'b00000010001011110000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N101.lt_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N101.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N98 [1] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [1] ),
            .I4 (),
            .ID ());
	// LUT = (~I2&~I3)|(I0&~I1&~I3)|(I0&~I1&~I2) ;
	// CARRY = (1'b0) ? CIN : ((~I2&~I3)|(I0&~I1&~I3)|(I0&~I1&~I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N101.lt_1  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N101.lt_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N101.co [2] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N101.co [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N100 [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N100 [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [3] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N101.lt_2  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N101.lt_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N101.co [4] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N101.co [2] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N100 [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N100 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [5] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N101.lt_3  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N101.lt_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N101.co [6] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N101.co [4] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N100 [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N100 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [7] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N101.lt_4  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N101.lt_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N101.co [8] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N101.co [6] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N100 [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N100 [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [9] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N101.lt_5  */ #(
            .INIT(32'b10100000111110100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N101.lt_5  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N101 ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N101.co [8] ),
            .I0 (),
            .I1 (),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N100 [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [10] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(CIN&~I3)|(CIN&I2) ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT1 /* \u_lcd_rgb_char/u_lcd_driver/N106_0_sum6_1  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_lcd_driver/N106_0_sum6_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/nb3 [6] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ));
	// LUT = ~I0 ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_0  */ #(
            .INIT(32'b11001100110011000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_0  (
            .COUT (_N645),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [1] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I1 ;
	// CARRY = (1'b0) ? CIN : (I1) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_1  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_1  (
            .COUT (_N646),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N106 [2] ),
            .CIN (_N645),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [2] ),
            .I2 (),
            .I3 (),
            .I4 (1'b1),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_2  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_2  (
            .COUT (_N647),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N106 [3] ),
            .CIN (_N646),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [3] ),
            .I2 (),
            .I3 (),
            .I4 (1'b1),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_3  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_3  (
            .COUT (_N648),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N106 [4] ),
            .CIN (_N647),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N98 [4] ),
            .I2 (),
            .I3 (),
            .I4 (1'b1),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_4  */ #(
            .INIT(32'b01011010011010011111000011000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_4  (
            .COUT (_N649),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N106 [5] ),
            .CIN (_N648),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N98 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [5] ),
            .ID ());
	// LUT = (~CIN&~I1&~I2&~I3)|(CIN&~I1&I2&~I3)|(CIN&~I2&I3)|(~CIN&I2&I3)|(CIN&I1&~I2)|(~CIN&I1&I2) ;
	// CARRY = ((~I1&~I2&~I3)|(I2&I3)|(I1&I2)) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_5  */ #(
            .INIT(32'b01101001011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_5  (
            .COUT (_N650),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N106 [6] ),
            .CIN (_N649),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N98 [6] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [6] ),
            .ID ());
	// LUT = ~I2^I1^CIN ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_6  */ #(
            .INIT(32'b01101001011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_6  (
            .COUT (_N651),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N106 [7] ),
            .CIN (_N650),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N98 [7] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [7] ),
            .ID ());
	// LUT = ~I2^I1^CIN ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_7  */ #(
            .INIT(32'b01101001011010011100001111000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_7  (
            .COUT (_N652),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N106 [8] ),
            .CIN (_N651),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N98 [8] ),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/N98 [8] ),
            .ID ());
	// LUT = ~I2^I1^CIN ;
	// CARRY = (~I2^I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_8  */ #(
            .INIT(32'b10101001101010010000001100000011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_8  (
            .COUT (_N653),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N106 [9] ),
            .CIN (_N652),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (~CIN&~I1&~I2)|(CIN&I2)|(CIN&I1) ;
	// CARRY = (~I1&~I2) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N106_2_9  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N106_2_9  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N106 [10] ),
            .CIN (_N653),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N107.lt_0  */ #(
            .INIT(32'b00000010001011110000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N107.lt_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N107.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [0] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N98 [1] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [1] ),
            .I4 (),
            .ID ());
	// LUT = (~I2&~I3)|(I0&~I1&~I3)|(I0&~I1&~I2) ;
	// CARRY = (1'b0) ? CIN : ((~I2&~I3)|(I0&~I1&~I3)|(I0&~I1&~I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N107.lt_1  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N107.lt_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N107.co [2] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N107.co [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N106 [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N106 [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [3] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N107.lt_2  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N107.lt_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N107.co [4] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N107.co [2] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N106 [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N106 [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [5] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N107.lt_3  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N107.lt_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N107.co [6] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N107.co [4] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N106 [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N106 [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [7] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N107.lt_4  */ #(
            .INIT(32'b00100000111100101001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N107.lt_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N107.co [8] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N107.co [6] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N106 [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N106 [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [9] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2) ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : ((I2&~I3)|(I0&~I1&~I3)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N107.lt_5  */ #(
            .INIT(32'b10100000111110100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N107.lt_5  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N107 ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N107.co [8] ),
            .I0 (),
            .I1 (),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N106 [10] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [10] ),
            .I4 (),
            .ID ());
	// LUT = (I2&~I3)|(CIN&~I3)|(CIN&I2) ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:227

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_driver/N116_5  */ #(
            .INIT(16'b0000010000000000))
        \u_lcd_rgb_char/u_lcd_driver/N116_5  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N116 ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N13 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N101 ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N107 ));
	// LUT = ~I0&I1&~I2&I3 ;

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_0  */ #(
            .INIT(32'b10101010101010100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I0 ;
	// CARRY = (1'b0) ? CIN : (I0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_1  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [1] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N124 [5] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [0] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [4] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_back [4] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_2  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [2] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N124 [6] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [1] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_3  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [3] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N124 [7] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [2] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_4  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [4] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N124 [8] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [3] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [10] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_disp [10] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_5  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_5  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [5] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N124 [9] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [4] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_6  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N124_1.fsub_6  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N124 [10] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N124_1.co [5] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_total [10] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_total [10] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N125.eq_0  */ #(
            .INIT(32'b00100100001001000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N125.eq_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N125.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [1] ),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = (~I0&I1&~I2)|(I0&~I1&I2) ;
	// CARRY = (1'b0) ? CIN : ((~I0&I1&~I2)|(I0&~I1&I2)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N125.eq_1  */ #(
            .INIT(32'b00000000000000001000100010001000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N125.eq_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N125.co [2] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N125.co [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [3] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = (I0&I1) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N125.eq_2  */ #(
            .INIT(32'b00000000000000000110000000000110), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N125.eq_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N125.co [4] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N125.co [2] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N124 [5] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((I0&~I1&~I2&~I3)|(~I0&I1&~I2&~I3)|(I0&~I1&I2&I3)|(~I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N125.eq_3  */ #(
            .INIT(32'b00000000000000001001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N125.eq_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N125.co [6] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N125.co [4] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N124 [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N124 [7] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N125.eq_4  */ #(
            .INIT(32'b00000000000000001001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N125.eq_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N125.co [8] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N125.co [6] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N124 [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N124 [9] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N125.eq_5  */ #(
            .INIT(32'b10100000000010100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N125.eq_5  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N125.co [8] ),
            .I0 (),
            .I1 (),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [10] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N124 [10] ),
            .I4 (),
            .ID ());
	// LUT = (CIN&~I2&~I3)|(CIN&I2&I3) ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:239

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_0  */ #(
            .INIT(32'b11001100110011000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_0  (
            .COUT (_N711),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [0] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I1 ;
	// CARRY = (1'b0) ? CIN : (I1) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_1  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_1  (
            .COUT (_N712),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [1] ),
            .CIN (_N711),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_2  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_2  (
            .COUT (_N713),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [2] ),
            .CIN (_N712),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_3  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_3  (
            .COUT (_N714),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [3] ),
            .CIN (_N713),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [3] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_4  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_4  (
            .COUT (_N715),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [4] ),
            .CIN (_N714),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_5  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_5  (
            .COUT (_N716),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [5] ),
            .CIN (_N715),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [5] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_6  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_6  (
            .COUT (_N717),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [6] ),
            .CIN (_N716),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_7  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_7  (
            .COUT (_N718),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [7] ),
            .CIN (_N717),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [7] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_8  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_8  (
            .COUT (_N719),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [8] ),
            .CIN (_N718),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_9  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_9  (
            .COUT (_N720),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [9] ),
            .CIN (_N719),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N132_1_10  */ #(
            .INIT(32'b00000110000001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N132_1_10  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [10] ),
            .CIN (_N720),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [10] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&~I2)|(~CIN&I1&~I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:242

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_0  */ #(
            .INIT(32'b00110011001100110000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [0] ),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = ~I1 ;
	// CARRY = (1'b0) ? CIN : (~I1) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_1  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [1] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [1] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [0] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb3 [6] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb3 [6] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_2  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [2] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [2] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [1] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [8] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_disp [8] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_3  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [3] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [3] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [2] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb3 [8] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb3 [8] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_4  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [4] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [4] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [3] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb3 [6] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/nb3 [6] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_5  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_5  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [5] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [5] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [4] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [10] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_disp [10] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_6  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_6  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [6] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [6] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [5] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_7  */ #(
            .INIT(32'b01010101010101011111111111111111), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_7  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [7] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [7] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [6] ),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~CIN ;
	// CARRY = (1'b1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_8  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_8  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [8] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [8] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [7] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_9  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_9  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [9] ),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [9] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [8] ),
            .I0 (),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_total [10] ),
            .I2 (),
            .I3 (),
            .I4 (\u_lcd_rgb_char/u_lcd_driver/h_total [10] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_10  */ #(
            .INIT(32'b01010101010101011111111111111111), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N144_1.fsub_10  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N144 [10] ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N144_1.co [9] ),
            .I0 (),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = ~CIN ;
	// CARRY = (1'b1) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N145.eq_0  */ #(
            .INIT(32'b10010000000010010000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N145.eq_0  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N145.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [0] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [1] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N144 [1] ),
            .I4 (),
            .ID ());
	// LUT = (~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3) ;
	// CARRY = (1'b0) ? CIN : ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N145.eq_1  */ #(
            .INIT(32'b00000000000000001001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N145.eq_1  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N145.co [2] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N145.co [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [2] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N144 [2] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [3] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N144 [3] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N145.eq_2  */ #(
            .INIT(32'b00000000000000001001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N145.eq_2  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N145.co [4] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N145.co [2] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [4] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N144 [4] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [5] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N144 [5] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N145.eq_3  */ #(
            .INIT(32'b00000000000000001001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N145.eq_3  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N145.co [6] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N145.co [4] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [6] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N144 [6] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [7] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N144 [7] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N145.eq_4  */ #(
            .INIT(32'b00000000000000001001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N145.eq_4  (
            .COUT (\u_lcd_rgb_char/u_lcd_driver/N145.co [8] ),
            .Z (),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N145.co [6] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [8] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N144 [8] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [9] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N144 [9] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT5CARRY /* \u_lcd_rgb_char/u_lcd_driver/N145.eq_5  */ #(
            .INIT(32'b10100000000010100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_lcd_rgb_char/u_lcd_driver/N145.eq_5  (
            .COUT (),
            .Z (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .CIN (\u_lcd_rgb_char/u_lcd_driver/N145.co [8] ),
            .I0 (),
            .I1 (),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [10] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/N144 [10] ),
            .I4 (),
            .ID ());
	// LUT = (CIN&~I2&~I3)|(CIN&I2&I3) ;
	// CARRY = (1'b0) ? CIN : (I4) ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:252

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[0]_1  */ #(
            .INIT(4'b0001))
        \u_lcd_rgb_char/u_lcd_driver/N153[0]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [0] ));
	// LUT = ~I0&~I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[1]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[1]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [1] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [1] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[2]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[2]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [2] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [2] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[3]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[3]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [3] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [3] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[4]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[4]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [4] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [4] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[5]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[5]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [5] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [5] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[6]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[6]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [6] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [6] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[7]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[7]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [7] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [7] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[8]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[8]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [8] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [8] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[9]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[9]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [9] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [9] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N153[10]_1  */ #(
            .INIT(4'b0100))
        \u_lcd_rgb_char/u_lcd_driver/N153[10]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N153 [10] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N145 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/N23 [10] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:255

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N178[0]_1  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_driver/N178[0]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N178 [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/nb1 [0] ));
	// LUT = I0&I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N180[0]_3  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_driver/N180[0]_3  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I1 (_N12225));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N180[1]_3  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_driver/N180[1]_3  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [1] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I1 (_N12226));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N180[2]_3  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_driver/N180[2]_3  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [2] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I1 (_N12227));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N180[3]_3  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_driver/N180[3]_3  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [3] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I1 (_N12228));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N180[4]_3  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_driver/N180[4]_3  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [4] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I1 (_N12229));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N180[5]_3  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_driver/N180[5]_3  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [5] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I1 (_N12230));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N180[6]_3  */ #(
            .INIT(4'b1000))
        \u_lcd_rgb_char/u_lcd_driver/N180[6]_3  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N180 [6] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N17 ),
            .I1 (_N12231));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/N182[0]_1  */ #(
            .INIT(4'b0001))
        \u_lcd_rgb_char/u_lcd_driver/N182[0]_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/N182 [0] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [0] ));
	// LUT = ~I0&~I1 ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_LUT3 /* \u_lcd_rgb_char/u_lcd_driver/N186_1  */ #(
            .INIT(8'b10101011))
        \u_lcd_rgb_char/u_lcd_driver/N186_1  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ),
            .I0 (\u_lcd_rgb_char/u_clk_div/N39 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ));
	// LUT = (~I1&~I2)|(I0) ;

    GTP_LUT1 /* \u_lcd_rgb_char/u_lcd_driver/N186_inv  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_lcd_driver/N186_inv  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_disp [8] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_back [2] ));
	// LUT = ~I0 ;

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/data_req  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/data_req_vname  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/data_req ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N116 ));
    // defparam \u_lcd_rgb_char/u_lcd_driver/data_req_vname .orig_name = \u_lcd_rgb_char/u_lcd_driver/data_req ;
	// ../../rtl/lcd_rgb_char/lcd_driver.v:224

    GTP_LUT2 /* \u_lcd_rgb_char/u_lcd_driver/h_back_or[1]  */ #(
            .INIT(4'b1110))
        \u_lcd_rgb_char/u_lcd_driver/h_back_or[1]  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_back [4] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT4 /* \u_lcd_rgb_char/u_lcd_driver/h_back_or[3]_2  */ #(
            .INIT(16'b1111101011111011))
        \u_lcd_rgb_char/u_lcd_driver/h_back_or[3]_2  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_disp [10] ),
            .I0 (\u_lcd_rgb_char/u_clk_div/N39 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_disp [9] ),
            .I2 (\u_lcd_rgb_char/u_lcd_driver/h_sync [1] ),
            .I3 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ));
	// LUT = (~I1&~I3)|(I2)|(I0) ;

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[0]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [0] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[1]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [1] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[2]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [2] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[3]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [3] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[4]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [4] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[5]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [5] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[6]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [6] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[7]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [7] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[8]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [8] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[9]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [9] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_LUT1 /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[10:0]_inv  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[10:0]_inv  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_cnt[1]_inv ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_cnt [1] ));
	// LUT = ~I0 ;

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/h_cnt[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/h_cnt[10]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/h_cnt [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N182 [10] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:235

    GTP_LUT1 /* \u_lcd_rgb_char/u_lcd_driver/h_total_inv  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_lcd_driver/h_total_inv  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/h_total [10] ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/h_back [1] ));
	// LUT = ~I0 ;

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/lcd_de  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/lcd_de  (
            .Q (nt_lcd_de),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/data_req ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:216

    GTP_LUT1 /* \u_lcd_rgb_char/u_lcd_driver/lcd_de_inv  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_lcd_driver/lcd_de_inv  (
            .Z (nt_lcd_de_inv),
            .I0 (nt_lcd_de));
	// LUT = ~I0 ;

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[0]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [0] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[1]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [1] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[2]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [2] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[3]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [3] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[4]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [4] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[5]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [5] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[6]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [6] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[7]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [7] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[8]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [8] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[9]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [9] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_xpos[10]  (
            .Q (\u_lcd_rgb_char/pixel_xpos_w [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N178 [10] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:130

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[0]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [0] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[1]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [1] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[2]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [2] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[3]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [3] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[4]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [4] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[5]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [5] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[6]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [6] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[7]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [7] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[8]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [8] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[9]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [9] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_LUT1 /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[10:0]_inv  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[10:0]_inv  (
            .Z (\u_lcd_rgb_char/pixel_ypos_w[0]_inv ),
            .I0 (\u_lcd_rgb_char/pixel_ypos_w [0] ));
	// LUT = ~I0 ;

    GTP_DFF_C /* \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/pixel_ypos[10]  (
            .Q (\u_lcd_rgb_char/pixel_ypos_w [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N180 [10] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:140

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[0]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [0] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[1]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [1] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[2]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [2] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[3]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [3] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[4]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [4] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[5]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [5] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[6]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [6] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[7]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [7] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[8]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [8] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[9]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [9] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_LUT1 /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[10:0]_inv  */ #(
            .INIT(2'b01))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[10:0]_inv  (
            .Z (\u_lcd_rgb_char/u_lcd_driver/v_cnt[0]_inv ),
            .I0 (\u_lcd_rgb_char/u_lcd_driver/v_cnt [0] ));
	// LUT = ~I0 ;

    GTP_DFF_CE /* \u_lcd_rgb_char/u_lcd_driver/v_cnt[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_lcd_driver/v_cnt[10]  (
            .Q (\u_lcd_rgb_char/u_lcd_driver/v_cnt [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_lcd_driver/N125 ),
            .CLK (nt_lcd_clk),
            .D (\u_lcd_rgb_char/u_lcd_driver/N153 [10] ));
	// ../../rtl/lcd_rgb_char/lcd_driver.v:247

    GTP_LUT3 /* \u_lcd_rgb_char/u_rd_id/N22_6[1]  */ #(
            .INIT(8'b00010110))
        \u_lcd_rgb_char/u_rd_id/N22_6[1]  (
            .Z (\u_lcd_rgb_char/u_rd_id/N22 [2] ),
            .I0 (_N0),
            .I1 (_N1),
            .I2 (_N2));
	// LUT = (I0&~I1&~I2)|(~I0&I1&~I2)|(~I0&~I1&I2) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_rd_id/N22_6[2]  */ #(
            .INIT(8'b00100100))
        \u_lcd_rgb_char/u_rd_id/N22_6[2]  (
            .Z (\u_lcd_rgb_char/u_rd_id/N22 [4] ),
            .I0 (_N0),
            .I1 (_N1),
            .I2 (_N2));
	// LUT = (~I0&I1&~I2)|(I0&~I1&I2) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_rd_id/N22_6[3]  */ #(
            .INIT(8'b00010010))
        \u_lcd_rgb_char/u_rd_id/N22_6[3]  (
            .Z (\u_lcd_rgb_char/u_rd_id/N22 [7] ),
            .I0 (_N0),
            .I1 (_N1),
            .I2 (_N2));
	// LUT = (I0&~I1&~I2)|(~I0&~I1&I2) ;

    GTP_LUT2 /* \u_lcd_rgb_char/u_rd_id/N22_6[4]  */ #(
            .INIT(4'b0001))
        \u_lcd_rgb_char/u_rd_id/N22_6[4]  (
            .Z (\u_lcd_rgb_char/u_rd_id/N22 [8] ),
            .I0 (_N1),
            .I1 (_N2));
	// LUT = ~I0&~I1 ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_rd_id/N22_6[5]  */ #(
            .INIT(8'b00110100))
        \u_lcd_rgb_char/u_rd_id/N22_6[5]  (
            .Z (\u_lcd_rgb_char/u_rd_id/N22 [12] ),
            .I0 (_N0),
            .I1 (_N1),
            .I2 (_N2));
	// LUT = (~I0&I1&~I2)|(~I1&I2) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_rd_id/N22_6[6]  */ #(
            .INIT(8'b00010100))
        \u_lcd_rgb_char/u_rd_id/N22_6[6]  (
            .Z (\u_lcd_rgb_char/u_rd_id/N22 [13] ),
            .I0 (_N0),
            .I1 (_N1),
            .I2 (_N2));
	// LUT = (~I0&I1&~I2)|(~I0&~I1&I2) ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_rd_id/N22_6[7]  */ #(
            .INIT(8'b00010111))
        \u_lcd_rgb_char/u_rd_id/N22_6[7]  (
            .Z (\u_lcd_rgb_char/u_rd_id/N22 [14] ),
            .I0 (_N0),
            .I1 (_N1),
            .I2 (_N2));
	// LUT = (~I1&~I2)|(~I0&~I2)|(~I0&~I1) ;

    GTP_INV \u_lcd_rgb_char/u_rd_id/N27_vname  (
            .Z (\u_lcd_rgb_char/u_rd_id/N27 ),
            .I (\u_lcd_rgb_char/u_rd_id/rd_flag ));
    // defparam \u_lcd_rgb_char/u_rd_id/N27_vname .orig_name = \u_lcd_rgb_char/u_rd_id/N27 ;

    GTP_LUT3 /* \u_lcd_rgb_char/u_rd_id/N31  */ #(
            .INIT(8'b00000001))
        \u_lcd_rgb_char/u_rd_id/N31_vname  (
            .Z (\u_lcd_rgb_char/u_rd_id/N31 ),
            .I0 (_N0),
            .I1 (_N1),
            .I2 (_N2));
    // defparam \u_lcd_rgb_char/u_rd_id/N31_vname .orig_name = \u_lcd_rgb_char/u_rd_id/N31 ;
	// LUT = ~I0&~I1&~I2 ;
	// ../../rtl/lcd_rgb_char/rd_id.v:43

    GTP_LUT3 /* \u_lcd_rgb_char/u_rd_id/N35  */ #(
            .INIT(8'b00100000))
        \u_lcd_rgb_char/u_rd_id/N35_vname  (
            .Z (\u_lcd_rgb_char/u_rd_id/N35 ),
            .I0 (_N0),
            .I1 (_N1),
            .I2 (_N2));
    // defparam \u_lcd_rgb_char/u_rd_id/N35_vname .orig_name = \u_lcd_rgb_char/u_rd_id/N35 ;
	// LUT = I0&~I1&I2 ;
	// ../../rtl/lcd_rgb_char/rd_id.v:47

    GTP_LUT2 /* \u_lcd_rgb_char/u_rd_id/N35_2  */ #(
            .INIT(4'b0001))
        \u_lcd_rgb_char/u_rd_id/N35_2  (
            .Z (\u_lcd_rgb_char/u_rd_id/N22 [1] ),
            .I0 (_N0),
            .I1 (_N2));
	// LUT = ~I0&~I1 ;

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[1]  (
            .Q (lcd_id[1]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N22 [1] ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[2]  (
            .Q (lcd_id[2]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N22 [2] ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[3]  (
            .Q (lcd_id[3]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N35 ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[4]  (
            .Q (lcd_id[4]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N22 [4] ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[6]  (
            .Q (lcd_id[6]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N31 ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[7]  (
            .Q (lcd_id[7]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N22 [7] ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[8]  (
            .Q (lcd_id[8]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N22 [8] ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[12]  (
            .Q (lcd_id[12]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N22 [12] ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[13]  (
            .Q (lcd_id[13]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N22 [13] ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/lcd_id[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/lcd_id[14]  (
            .Q (lcd_id[14]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (\u_lcd_rgb_char/u_rd_id/N22 [14] ));
	// ../../rtl/lcd_rgb_char/rd_id.v:34

    GTP_DFF_CE /* \u_lcd_rgb_char/u_rd_id/rd_flag  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_lcd_rgb_char/u_rd_id/rd_flag_vname  (
            .Q (\u_lcd_rgb_char/u_rd_id/rd_flag ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_lcd_rgb_char/u_rd_id/N27 ),
            .CLK (nt_sys_clk),
            .D (1'b1));
    // defparam \u_lcd_rgb_char/u_rd_id/rd_flag_vname .orig_name = \u_lcd_rgb_char/u_rd_id/rd_flag ;
	// ../../rtl/lcd_rgb_char/rd_id.v:34

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="J3", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_IOBUF /* \u_touch_top.u_i2c_dri.sda_tri  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"), 
            .TERM_DDR("ON"))
        \u_touch_top.u_i2c_dri.sda_tri  (
            .IO (touch_sda),
            .O (_N3),
            .I (\u_touch_top/u_i2c_dri/sda_out ),
            .T (\u_touch_top/u_i2c_dri/sda_dir_inv ));
	// ../../rtl/top_lcd_touch.v:23

(* PAP_IO_DIRECTION="INOUT", PAP_IO_LOC="F3", PAP_IO_VCCIO="3.3", PAP_IO_STANDARD="LVCMOS33", PAP_IO_DRIVE="8", PAP_IO_PULLUP="TRUE", PAP_IO_SLEW="SLOW" *)    GTP_OUTBUFT /* \u_touch_top.u_touch_dri.touch_int_tri  */ #(
            .IOSTANDARD("DEFAULT"), 
            .SLEW_RATE("SLOW"), 
            .DRIVE_STRENGTH("8"))
        \u_touch_top.u_touch_dri.touch_int_tri  (
            .O (touch_int),
            .I (\u_touch_top/u_touch_dri/touch_int_out ),
            .T (\u_touch_top/u_touch_dri/touch_int_dir_inv ));
	// ../../rtl/top_lcd_touch.v:25

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N2.eq_0  */ #(
            .INIT(32'b10010000000010010000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N2.eq_0  (
            .COUT (\u_touch_top/u_i2c_dri/N2.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_touch_top/reg_num [0] ),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [0] ),
            .I2 (\u_touch_top/reg_num [1] ),
            .I3 (\u_touch_top/u_i2c_dri/reg_cnt [1] ),
            .I4 (),
            .ID ());
	// LUT = (~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3) ;
	// CARRY = (1'b0) ? CIN : ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ;
	// ../../rtl/touch/i2c_dri.v:83

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N2.eq_1  */ #(
            .INIT(32'b00000000000000000000100100001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N2.eq_1  (
            .COUT (\u_touch_top/u_i2c_dri/N2.co [2] ),
            .Z (),
            .CIN (\u_touch_top/u_i2c_dri/N2.co [0] ),
            .I0 (\u_touch_top/reg_num [2] ),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/reg_cnt [3] ),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2)|(I0&I1&~I2)) ? CIN : (1'b0) ;
	// ../../rtl/touch/i2c_dri.v:83

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N2.eq_2  */ #(
            .INIT(32'b00000000000000000000000000000001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N2.eq_2  (
            .COUT (\u_touch_top/u_i2c_dri/reg_done ),
            .Z (),
            .CIN (\u_touch_top/u_i2c_dri/N2.co [2] ),
            .I0 (\u_touch_top/u_i2c_dri/reg_cnt [4] ),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [5] ),
            .I2 (\u_touch_top/u_i2c_dri/reg_cnt [6] ),
            .I3 (\u_touch_top/u_i2c_dri/reg_cnt [7] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = (~I0&~I1&~I2&~I3) ? CIN : (1'b0) ;
	// ../../rtl/touch/i2c_dri.v:83

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N12_1_0  */ #(
            .INIT(32'b11001100110011000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N12_1_0  (
            .COUT (_N722),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [0] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I1 ;
	// CARRY = (1'b0) ? CIN : (I1) ;
	// ../../rtl/touch/i2c_dri.v:96

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N12_1_1  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N12_1_1  (
            .COUT (_N723),
            .Z (\u_touch_top/u_i2c_dri/N12 [1] ),
            .CIN (_N722),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [1] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:96

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N12_1_2  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N12_1_2  (
            .COUT (_N724),
            .Z (\u_touch_top/u_i2c_dri/N12 [2] ),
            .CIN (_N723),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [2] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:96

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N12_1_3  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N12_1_3  (
            .COUT (_N725),
            .Z (\u_touch_top/u_i2c_dri/N12 [3] ),
            .CIN (_N724),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [3] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:96

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N12_1_4  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N12_1_4  (
            .COUT (_N726),
            .Z (\u_touch_top/u_i2c_dri/N811 [4] ),
            .CIN (_N725),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [4] ),
            .I2 (\u_touch_top/u_i2c_dri/N582_inv ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:96

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N12_1_5  */ #(
            .INIT(32'b00100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N12_1_5  (
            .COUT (),
            .Z (\u_touch_top/u_i2c_dri/N811 [5] ),
            .CIN (_N726),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [5] ),
            .I2 (\u_touch_top/u_i2c_dri/clk_cnt [0] ),
            .I3 (_N12050),
            .I4 (1'b0),
            .ID ());
	// LUT = (~CIN&I1&~I3)|(~CIN&I1&~I2)|(CIN&~I1) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:96

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N20_1_0  */ #(
            .INIT(32'b11001100110011000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N20_1_0  (
            .COUT (_N682),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [0] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I1 ;
	// CARRY = (1'b0) ? CIN : (I1) ;
	// ../../rtl/touch/i2c_dri.v:104

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N20_1_1  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N20_1_1  (
            .COUT (_N683),
            .Z (\u_touch_top/u_i2c_dri/N815 [1] ),
            .CIN (_N682),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [1] ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:104

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N20_1_2  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N20_1_2  (
            .COUT (_N684),
            .Z (\u_touch_top/u_i2c_dri/N815 [2] ),
            .CIN (_N683),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [2] ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:104

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N20_1_3  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N20_1_3  (
            .COUT (_N685),
            .Z (\u_touch_top/u_i2c_dri/N815 [3] ),
            .CIN (_N684),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [3] ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:104

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N20_1_4  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N20_1_4  (
            .COUT (_N686),
            .Z (\u_touch_top/u_i2c_dri/N815 [4] ),
            .CIN (_N685),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [4] ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:104

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N20_1_5  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N20_1_5  (
            .COUT (_N687),
            .Z (\u_touch_top/u_i2c_dri/N815 [5] ),
            .CIN (_N686),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [5] ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:104

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N20_1_6  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N20_1_6  (
            .COUT (_N688),
            .Z (\u_touch_top/u_i2c_dri/N815 [6] ),
            .CIN (_N687),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [6] ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:104

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N20_1_7  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N20_1_7  (
            .COUT (),
            .Z (\u_touch_top/u_i2c_dri/N815 [7] ),
            .CIN (_N688),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [7] ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:104

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N97_1_0  */ #(
            .INIT(32'b11001100110011000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N97_1_0  (
            .COUT (_N675),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I1 ;
	// CARRY = (1'b0) ? CIN : (I1) ;
	// ../../rtl/touch/i2c_dri.v:226

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N97_1_1  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N97_1_1  (
            .COUT (_N676),
            .Z (\u_touch_top/u_i2c_dri/N97 [1] ),
            .CIN (_N675),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:226

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N97_1_2  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N97_1_2  (
            .COUT (_N677),
            .Z (\u_touch_top/u_i2c_dri/N97 [2] ),
            .CIN (_N676),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:226

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N97_1_3  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N97_1_3  (
            .COUT (_N678),
            .Z (\u_touch_top/u_i2c_dri/N97 [3] ),
            .CIN (_N677),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:226

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N97_1_4  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N97_1_4  (
            .COUT (_N679),
            .Z (\u_touch_top/u_i2c_dri/N97 [4] ),
            .CIN (_N678),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:226

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N97_1_5  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N97_1_5  (
            .COUT (_N680),
            .Z (\u_touch_top/u_i2c_dri/N97 [5] ),
            .CIN (_N679),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:226

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N97_1_6  */ #(
            .INIT(32'b01100110011001101100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N97_1_6  (
            .COUT (),
            .Z (\u_touch_top/u_i2c_dri/N97 [6] ),
            .CIN (_N680),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/cnt [6] ),
            .I2 (),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = I1^CIN ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:226

    GTP_ROM32X1 /* \u_touch_top/u_i2c_dri/N171_2  */ #(
            .INIT(32'b00000000000000000000010000000000))
        \u_touch_top/u_i2c_dri/N171_2  (
            .Z (_N728),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [4] ));

    GTP_ROM32X1 /* \u_touch_top/u_i2c_dri/N237_2  */ #(
            .INIT(32'b00000000000000000000000001000000))
        \u_touch_top/u_i2c_dri/N237_2  (
            .Z (_N729),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [4] ));

    GTP_ROM32X1 /* \u_touch_top/u_i2c_dri/N369_2  */ #(
            .INIT(32'b00000000000000000000000000000001))
        \u_touch_top/u_i2c_dri/N369_2  (
            .Z (_N730),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [4] ));

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N475_1.fsub_0  */ #(
            .INIT(32'b10101010101010100000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N475_1.fsub_0  (
            .COUT (\u_touch_top/u_i2c_dri/N475_1.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_touch_top/u_i2c_dri/reg_cnt [0] ),
            .I1 (),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I0 ;
	// CARRY = (1'b0) ? CIN : (I0) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N475_1.fsub_1  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N475_1.fsub_1  (
            .COUT (\u_touch_top/u_i2c_dri/N475_1.co [1] ),
            .Z (\u_touch_top/u_i2c_dri/N475 [1] ),
            .CIN (\u_touch_top/u_i2c_dri/N475_1.co [0] ),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [1] ),
            .I2 (),
            .I3 (),
            .I4 (\u_touch_top/u_i2c_dri/reg_cnt [1] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N475_1.fsub_2  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N475_1.fsub_2  (
            .COUT (\u_touch_top/u_i2c_dri/N475_1.co [2] ),
            .Z (\u_touch_top/u_i2c_dri/N475 [2] ),
            .CIN (\u_touch_top/u_i2c_dri/N475_1.co [1] ),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [2] ),
            .I2 (),
            .I3 (),
            .I4 (\u_touch_top/u_i2c_dri/reg_cnt [2] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N475_1.fsub_3  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N475_1.fsub_3  (
            .COUT (\u_touch_top/u_i2c_dri/N475_1.co [3] ),
            .Z (\u_touch_top/u_i2c_dri/N475 [3] ),
            .CIN (\u_touch_top/u_i2c_dri/N475_1.co [2] ),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [3] ),
            .I2 (),
            .I3 (),
            .I4 (\u_touch_top/u_i2c_dri/reg_cnt [3] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N475_1.fsub_4  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N475_1.fsub_4  (
            .COUT (\u_touch_top/u_i2c_dri/N475_1.co [4] ),
            .Z (\u_touch_top/u_i2c_dri/N475 [4] ),
            .CIN (\u_touch_top/u_i2c_dri/N475_1.co [3] ),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [4] ),
            .I2 (),
            .I3 (),
            .I4 (\u_touch_top/u_i2c_dri/reg_cnt [4] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N475_1.fsub_5  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N475_1.fsub_5  (
            .COUT (\u_touch_top/u_i2c_dri/N475_1.co [5] ),
            .Z (\u_touch_top/u_i2c_dri/N475 [5] ),
            .CIN (\u_touch_top/u_i2c_dri/N475_1.co [4] ),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [5] ),
            .I2 (),
            .I3 (),
            .I4 (\u_touch_top/u_i2c_dri/reg_cnt [5] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N475_1.fsub_6  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N475_1.fsub_6  (
            .COUT (\u_touch_top/u_i2c_dri/N475_1.co [6] ),
            .Z (\u_touch_top/u_i2c_dri/N475 [6] ),
            .CIN (\u_touch_top/u_i2c_dri/N475_1.co [5] ),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [6] ),
            .I2 (),
            .I3 (),
            .I4 (\u_touch_top/u_i2c_dri/reg_cnt [6] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N475_1.fsub_7  */ #(
            .INIT(32'b10011001100110010011001100110011), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N475_1.fsub_7  (
            .COUT (),
            .Z (\u_touch_top/u_i2c_dri/N475 [7] ),
            .CIN (\u_touch_top/u_i2c_dri/N475_1.co [6] ),
            .I0 (),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [7] ),
            .I2 (),
            .I3 (),
            .I4 (\u_touch_top/u_i2c_dri/reg_cnt [7] ),
            .ID ());
	// LUT = ~I1^CIN ;
	// CARRY = (~I1) ? CIN : (I4) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N476.eq_0  */ #(
            .INIT(32'b00000000000000000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N476.eq_0  (
            .COUT (\u_touch_top/u_i2c_dri/N476.co [0] ),
            .Z (),
            .CIN (),
            .I0 (\u_touch_top/u_i2c_dri/reg_cnt [0] ),
            .I1 (),
            .I2 (\u_touch_top/u_i2c_dri/reg_cnt [1] ),
            .I3 (\u_touch_top/u_i2c_dri/N475 [1] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = (1'b0) ? CIN : (1'b0) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N476.eq_1  */ #(
            .INIT(32'b00000000000000001001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N476.eq_1  (
            .COUT (\u_touch_top/u_i2c_dri/N476.co [2] ),
            .Z (),
            .CIN (\u_touch_top/u_i2c_dri/N476.co [0] ),
            .I0 (\u_touch_top/u_i2c_dri/reg_cnt [2] ),
            .I1 (\u_touch_top/u_i2c_dri/N475 [2] ),
            .I2 (\u_touch_top/u_i2c_dri/reg_cnt [3] ),
            .I3 (\u_touch_top/u_i2c_dri/N475 [3] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N476.eq_2  */ #(
            .INIT(32'b00000000000000001001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N476.eq_2  (
            .COUT (\u_touch_top/u_i2c_dri/N476.co [4] ),
            .Z (),
            .CIN (\u_touch_top/u_i2c_dri/N476.co [2] ),
            .I0 (\u_touch_top/u_i2c_dri/reg_cnt [4] ),
            .I1 (\u_touch_top/u_i2c_dri/N475 [4] ),
            .I2 (\u_touch_top/u_i2c_dri/reg_cnt [5] ),
            .I3 (\u_touch_top/u_i2c_dri/N475 [5] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_LUT5CARRY /* \u_touch_top/u_i2c_dri/N476.eq_3  */ #(
            .INIT(32'b00000000000000001001000000001001), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_i2c_dri/N476.eq_3  (
            .COUT (\u_touch_top/u_i2c_dri/N476 ),
            .Z (),
            .CIN (\u_touch_top/u_i2c_dri/N476.co [4] ),
            .I0 (\u_touch_top/u_i2c_dri/reg_cnt [6] ),
            .I1 (\u_touch_top/u_i2c_dri/N475 [6] ),
            .I2 (\u_touch_top/u_i2c_dri/reg_cnt [7] ),
            .I3 (\u_touch_top/u_i2c_dri/N475 [7] ),
            .I4 (),
            .ID ());
	// LUT = 1'b0 ;
	// CARRY = ((~I0&~I1&~I2&~I3)|(I0&I1&~I2&~I3)|(~I0&~I1&I2&I3)|(I0&I1&I2&I3)) ? CIN : (1'b0) ;
	// ../../rtl/touch/i2c_dri.v:517

    GTP_ROM32X1 /* \u_touch_top/u_i2c_dri/N514_2  */ #(
            .INIT(32'b00000000000000000000000000000010))
        \u_touch_top/u_i2c_dri/N514_2  (
            .Z (_N731),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [4] ));

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N552_2  */ #(
            .INIT(16'b1111111111111110))
        \u_touch_top/u_i2c_dri/N552_2  (
            .Z (\u_touch_top/u_i2c_dri/_N42 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT3 /* \u_touch_top/u_i2c_dri/N552_4  */ #(
            .INIT(8'b00110010))
        \u_touch_top/u_i2c_dri/N552_4  (
            .Z (_N784),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_i2c_dri/N637 ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ));
	// LUT = (~I1&I2)|(I0&~I1) ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N552_6  */ #(
            .INIT(16'b1000000000000000))
        \u_touch_top/u_i2c_dri/N552_6  (
            .Z (_N785),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/_N42 ),
            .I3 (_N10567));
	// LUT = I0&I1&I2&I3 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N552_14_and[0][2]  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_i2c_dri/N552_14_and[0][2]  (
            .Z (\u_touch_top/u_i2c_dri/N552 [0] ),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (_N791));
	// LUT = ~I0&I1 ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N552_14_and[3][2]  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_i2c_dri/N552_14_and[3][2]  (
            .Z (\u_touch_top/u_i2c_dri/N552 [3] ),
            .I0 (\u_touch_top/u_i2c_dri/N97 [3] ),
            .I1 (_N791));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N552_14_and[5][2]  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_i2c_dri/N552_14_and[5][2]  (
            .Z (\u_touch_top/u_i2c_dri/N552 [5] ),
            .I0 (\u_touch_top/u_i2c_dri/N97 [5] ),
            .I1 (_N791));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N552_14_or[1]_1  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_i2c_dri/N552_14_or[1]_1  (
            .Z (\u_touch_top/u_i2c_dri/N552 [1] ),
            .I0 (\u_touch_top/u_i2c_dri/N97 [1] ),
            .I1 (_N10233));
	// LUT = I0&I1 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N552_14_or[1]_2  */ #(
            .INIT(32'b11111111111111111111111111001000))
        \u_touch_top/u_i2c_dri/N552_14_or[1]_2  (
            .Z (_N10233),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_i2c_dri/N637 ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I3 (_N785),
            .I4 (_N791));
	// LUT = (I4)|(I3)|(I1&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N552_14_or[2]_1  */ #(
            .INIT(32'b10101000101000001010000010100000))
        \u_touch_top/u_i2c_dri/N552_14_or[2]_1  (
            .Z (\u_touch_top/u_i2c_dri/N552 [2] ),
            .I0 (\u_touch_top/u_i2c_dri/N97 [2] ),
            .I1 (\u_touch_top/u_i2c_dri/_N42 ),
            .I2 (_N791),
            .I3 (_N10547),
            .I4 (_N10567));
	// LUT = (I0&I1&I3&I4)|(I0&I2) ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N552_14_or[4]_1  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_i2c_dri/N552_14_or[4]_1  (
            .Z (\u_touch_top/u_i2c_dri/N552 [4] ),
            .I0 (\u_touch_top/u_i2c_dri/N97 [4] ),
            .I1 (_N10233));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N552_14_or[6]_1  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_i2c_dri/N552_14_or[6]_1  (
            .Z (\u_touch_top/u_i2c_dri/N552 [6] ),
            .I0 (\u_touch_top/u_i2c_dri/N97 [6] ),
            .I1 (_N10233));
	// LUT = I0&I1 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N552_17_2  */ #(
            .INIT(32'b11111111011100001111111111110000))
        \u_touch_top/u_i2c_dri/N552_17_2  (
            .Z (_N11998),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/_N42 ),
            .I3 (_N784),
            .I4 (_N10567));
	// LUT = (I2&~I4)|(I3)|(~I1&I2)|(~I0&I2) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N552_17_3  */ #(
            .INIT(32'b11111111111111111000101010101010))
        \u_touch_top/u_i2c_dri/N552_17_3  (
            .Z (_N791),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [7] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N10568),
            .I4 (_N11998));
	// LUT = (I4)|(I0&~I3)|(I0&~I2)|(I0&I1) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N557_2_or[0]_1  */ #(
            .INIT(32'b11101010110000001100000011000000))
        \u_touch_top/u_i2c_dri/N557_2_or[0]_1  (
            .Z (\u_touch_top/u_i2c_dri/N557 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [7] ),
            .I1 (_N10361),
            .I2 (_N10483),
            .I3 (_N10547),
            .I4 (_N10569));
	// LUT = (I0&I3&I4)|(I1&I2) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N557_2_or[0]_5  */ #(
            .INIT(32'b11111110111100001110111000000000))
        \u_touch_top/u_i2c_dri/N557_2_or[0]_5  (
            .Z (_N10361),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I2 (\u_touch_top/u_i2c_dri/_N42 ),
            .I3 (_N728),
            .I4 (_N729));
	// LUT = (I2&I4)|(I1&I3)|(I0&I3) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N558_1_or[0]_1  */ #(
            .INIT(32'b11101010110000000000000000000000))
        \u_touch_top/u_i2c_dri/N558_1_or[0]_1  (
            .Z (\u_touch_top/u_i2c_dri/N558 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I2 (_N730),
            .I3 (_N731),
            .I4 (_N10483));
	// LUT = (I0&I3&I4)|(I1&I2&I4) ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N558_1_or[0]_6  */ #(
            .INIT(4'b0010))
        \u_touch_top/u_i2c_dri/N558_1_or[0]_6  (
            .Z (_N10483),
            .I0 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [6] ));
	// LUT = I0&~I1 ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N558_1_or[0]_7  */ #(
            .INIT(4'b0010))
        \u_touch_top/u_i2c_dri/N558_1_or[0]_7  (
            .Z (_N10545),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ));
	// LUT = I0&~I1 ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N558_1_or[0]_8  */ #(
            .INIT(4'b0001))
        \u_touch_top/u_i2c_dri/N558_1_or[0]_8  (
            .Z (_N10546),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ));
	// LUT = ~I0&~I1 ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N558_1_or[0]_9  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_i2c_dri/N558_1_or[0]_9  (
            .Z (_N10547),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ));
	// LUT = I0&I1 ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N558_1_or[0]_10  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_i2c_dri/N558_1_or[0]_10  (
            .Z (_N10548),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ));
	// LUT = ~I0&I1 ;

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N582_5  */ #(
            .INIT(16'b0000000100000000))
        \u_touch_top/u_i2c_dri/N582_5  (
            .Z (_N12050),
            .I0 (\u_touch_top/u_i2c_dri/clk_cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/clk_cnt [3] ),
            .I3 (\u_touch_top/u_i2c_dri/clk_cnt [4] ));
	// LUT = ~I0&~I1&~I2&I3 ;

    GTP_LUT3 /* \u_touch_top/u_i2c_dri/N582_inv  */ #(
            .INIT(8'b01111111))
        \u_touch_top/u_i2c_dri/N582_inv_vname  (
            .Z (\u_touch_top/u_i2c_dri/N582_inv ),
            .I0 (\u_touch_top/u_i2c_dri/clk_cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [5] ),
            .I2 (_N12050));
    // defparam \u_touch_top/u_i2c_dri/N582_inv_vname .orig_name = \u_touch_top/u_i2c_dri/N582_inv ;
	// LUT = (~I2)|(~I1)|(~I0) ;

    GTP_LUT3 /* \u_touch_top/u_i2c_dri/N607  */ #(
            .INIT(8'b00100000))
        \u_touch_top/u_i2c_dri/N607_vname  (
            .Z (\u_touch_top/u_i2c_dri/N607 ),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (_N10569));
    // defparam \u_touch_top/u_i2c_dri/N607_vname .orig_name = \u_touch_top/u_i2c_dri/N607 ;
	// LUT = I0&~I1&I2 ;
	// ../../rtl/touch/i2c_dri.v:242

    GTP_LUT3 /* \u_touch_top/u_i2c_dri/N607_1  */ #(
            .INIT(8'b00000001))
        \u_touch_top/u_i2c_dri/N607_1  (
            .Z (_N10539),
            .I0 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [6] ));
	// LUT = ~I0&~I1&~I2 ;

    GTP_LUT3 /* \u_touch_top/u_i2c_dri/N607_2  */ #(
            .INIT(8'b00000010))
        \u_touch_top/u_i2c_dri/N607_2  (
            .Z (_N10540),
            .I0 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [6] ));
	// LUT = I0&~I1&~I2 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N607_3  */ #(
            .INIT(32'b00000000000000000000000100000000))
        \u_touch_top/u_i2c_dri/N607_3  (
            .Z (_N10566),
            .I0 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [6] ));
	// LUT = ~I0&~I1&~I2&I3&~I4 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N607_4  */ #(
            .INIT(32'b00000000000000000000001000000000))
        \u_touch_top/u_i2c_dri/N607_4  (
            .Z (_N10567),
            .I0 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [6] ));
	// LUT = I0&~I1&~I2&I3&~I4 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N608_1  */ #(
            .INIT(32'b00000000000000000000000000000010))
        \u_touch_top/u_i2c_dri/N608_1  (
            .Z (_N10568),
            .I0 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [6] ));
	// LUT = I0&~I1&~I2&~I3&~I4 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N614_1  */ #(
            .INIT(32'b00000000000000000000000000000001))
        \u_touch_top/u_i2c_dri/N614_1  (
            .Z (_N10569),
            .I0 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [6] ));
	// LUT = ~I0&~I1&~I2&~I3&~I4 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N615_1  */ #(
            .INIT(32'b00000000000000000000000000010000))
        \u_touch_top/u_i2c_dri/N615_1  (
            .Z (_N10570),
            .I0 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [6] ));
	// LUT = ~I0&~I1&I2&~I3&~I4 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N621_1  */ #(
            .INIT(32'b00000000000000000000000001000000))
        \u_touch_top/u_i2c_dri/N621_1  (
            .Z (_N10571),
            .I0 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [5] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [6] ));
	// LUT = ~I0&I1&I2&~I3&~I4 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N637_7  */ #(
            .INIT(32'b00001000000000000000000000000000))
        \u_touch_top/u_i2c_dri/N637_7  (
            .Z (\u_touch_top/u_i2c_dri/N637 ),
            .I0 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (_N10483),
            .I4 (_N10545));
	// LUT = I0&I1&~I2&I3&I4 ;

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N811[0]  */ #(
            .INIT(16'b0010101010101010))
        \u_touch_top/u_i2c_dri/N811[0]  (
            .Z (\u_touch_top/u_i2c_dri/N811 [1] ),
            .I0 (\u_touch_top/u_i2c_dri/N12 [1] ),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/clk_cnt [5] ),
            .I3 (_N12050));
	// LUT = (I0&~I3)|(I0&~I2)|(I0&~I1) ;
	// ../../rtl/touch/i2c_dri.v:86

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N814  */ #(
            .INIT(4'b1110))
        \u_touch_top/u_i2c_dri/N814_vname  (
            .Z (\u_touch_top/u_i2c_dri/N814 ),
            .I0 (\u_touch_top/i2c_done ),
            .I1 (\u_touch_top/once_byte_done ));
    // defparam \u_touch_top/u_i2c_dri/N814_vname .orig_name = \u_touch_top/u_i2c_dri/N814 ;
	// LUT = (I1)|(I0) ;
	// ../../rtl/touch/i2c_dri.v:100

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N815[0]_1  */ #(
            .INIT(4'b0010))
        \u_touch_top/u_i2c_dri/N815[0]_1  (
            .Z (\u_touch_top/u_i2c_dri/N815 [0] ),
            .I0 (\u_touch_top/once_byte_done ),
            .I1 (\u_touch_top/u_i2c_dri/reg_cnt [0] ));
	// LUT = I0&~I1 ;
	// ../../rtl/touch/i2c_dri.v:100

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1180  */ #(
            .INIT(32'b11111111111111111010101010000000))
        \u_touch_top/u_i2c_dri/N1180_vname  (
            .Z (\u_touch_top/u_i2c_dri/N1180 ),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (_N10567),
            .I3 (_N10568),
            .I4 (_N11014_3));
    // defparam \u_touch_top/u_i2c_dri/N1180_vname .orig_name = \u_touch_top/u_i2c_dri/N1180 ;
	// LUT = (I4)|(I0&I3)|(I0&I1&I2) ;
	// ../../rtl/touch/i2c_dri.v:474

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1180_28  */ #(
            .INIT(32'b10101010101000000000000000000000))
        \u_touch_top/u_i2c_dri/N1180_28  (
            .Z (_N11014_3),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I4 (_N10540));
	// LUT = (I0&I3&I4)|(I0&I2&I4) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1181_11  */ #(
            .INIT(32'b00000010101010000000000000000000))
        \u_touch_top/u_i2c_dri/N1181_11  (
            .Z (_N12216),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I4 (_N10539));
	// LUT = (I0&I2&~I3&I4)|(I0&I1&~I3&I4)|(I0&~I1&~I2&I3&I4) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1181_13  */ #(
            .INIT(32'b11111111110010001111111111001000))
        \u_touch_top/u_i2c_dri/N1181_13  (
            .Z (_N10592),
            .I0 (_N10570),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (_N10571),
            .I3 (_N12216),
            .I4 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .ID (_N10566));
	// LUT = (ID&I1&~I4)|(I0&I1&I4)|(I3)|(I1&I2) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1185_5  */ #(
            .INIT(32'b11111111111111101111111111101100))
        \u_touch_top/u_i2c_dri/N1185_5  (
            .Z (\u_touch_top/u_i2c_dri/N1185 ),
            .I0 (_N10567),
            .I1 (\u_touch_top/u_i2c_dri/N637 ),
            .I2 (_N10568),
            .I3 (_N11014_3),
            .I4 (_N10545),
            .ID (_N10547));
	// LUT = (I2&I4)|(I0&I4)|(I3)|(ID&I2)|(I1) ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N1222  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_i2c_dri/N1222_vname  (
            .Z (\u_touch_top/u_i2c_dri/N1222 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/N1180 ));
    // defparam \u_touch_top/u_i2c_dri/N1222_vname .orig_name = \u_touch_top/u_i2c_dri/N1222 ;
	// LUT = I0&I1 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1227_1_2  */ #(
            .INIT(32'b11111111111010101010101010000000))
        \u_touch_top/u_i2c_dri/N1227_1_2  (
            .Z (_N12219),
            .I0 (\u_touch_top/u_i2c_dri/N607 ),
            .I1 (_N10547),
            .I2 (_N10566),
            .I3 (_N10592),
            .I4 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .ID (\u_touch_top/u_i2c_dri/cur_state_reg [1] ));
	// LUT = (I3&I4)|(I1&I2&I4)|(I0&I4)|(ID&I3)|(ID&I1&I2) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1227_1_3  */ #(
            .INIT(32'b10101010111010100000000010000000))
        \u_touch_top/u_i2c_dri/N1227_1_3  (
            .Z (_N12220),
            .I0 (_N10592),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (_N10569),
            .I3 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I4 (\u_touch_top/u_i2c_dri/_N42 ),
            .ID (\u_touch_top/u_i2c_dri/cur_state_reg [7] ));
	// LUT = (I1&I2&~I3&I4)|(I0&I4)|(ID&I1&I2&~I3) ;

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N1227_1_6  */ #(
            .INIT(16'b1111111111111110))
        \u_touch_top/u_i2c_dri/N1227_1_6  (
            .Z (\u_touch_top/u_i2c_dri/N1227 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [0] ),
            .I1 (\u_touch_top/u_i2c_dri/N1230 ),
            .I2 (_N12219),
            .I3 (_N12220));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1227_10  */ #(
            .INIT(32'b00110000001000000010000000100000))
        \u_touch_top/u_i2c_dri/N1227_10  (
            .Z (_N12010),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (_N10566),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .ID (_N11792_3));
	// LUT = (ID&~I1&I2&~I4)|(~I1&I2&I3&I4)|(I0&~I1&I2&I4) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1227_14  */ #(
            .INIT(32'b11111111111111110000001000000000))
        \u_touch_top/u_i2c_dri/N1227_14  (
            .Z (\u_touch_top/u_i2c_dri/N2082 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N10569),
            .I4 (_N12010));
	// LUT = (I4)|(I0&~I1&~I2&I3) ;

    GTP_LUT3 /* \u_touch_top/u_i2c_dri/N1230_8  */ #(
            .INIT(8'b11111110))
        \u_touch_top/u_i2c_dri/N1230_8  (
            .Z (_N11792_3),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ));
	// LUT = (I2)|(I1)|(I0) ;

    GTP_LUT1 /* \u_touch_top/u_i2c_dri/N1232  */ #(
            .INIT(2'b01))
        \u_touch_top/u_i2c_dri/N1232_vname  (
            .Z (\u_touch_top/u_i2c_dri/N1232 ),
            .I0 (\u_touch_top/u_i2c_dri/N1230 ));
    // defparam \u_touch_top/u_i2c_dri/N1232_vname .orig_name = \u_touch_top/u_i2c_dri/N1232 ;
	// LUT = ~I0 ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1596_9  */ #(
            .INIT(32'b11111111111101000000000000000000))
        \u_touch_top/u_i2c_dri/N1596_9  (
            .Z (_N11426_3),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I4 (_N10539));
	// LUT = (I3&I4)|(I2&I4)|(~I0&I1&I4) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1600  */ #(
            .INIT(32'b01010101010101010001000100010000))
        \u_touch_top/u_i2c_dri/N1600_vname  (
            .Z (\u_touch_top/u_i2c_dri/N1600 ),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (_N10566),
            .I3 (_N10569),
            .I4 (_N11426_3));
    // defparam \u_touch_top/u_i2c_dri/N1600_vname .orig_name = \u_touch_top/u_i2c_dri/N1600 ;
	// LUT = (~I0&I4)|(~I0&~I1&I3)|(~I0&~I1&I2) ;
	// ../../rtl/touch/i2c_dri.v:378

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1668_1_4  */ #(
            .INIT(32'b11111101111111111111110011111111))
        \u_touch_top/u_i2c_dri/N1668_1_4  (
            .Z (\u_touch_top/u_i2c_dri/N1668 ),
            .I0 (\u_touch_top/u_i2c_dri/N1600 ),
            .I1 (_N10344),
            .I2 (_N10345),
            .I3 (_N10992_1),
            .I4 (_N11792_3));
	// LUT = (~I0&I4)|(~I3)|(I2)|(I1) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1668_1_7  */ #(
            .INIT(32'b10001010110011110000000010001111))
        \u_touch_top/u_i2c_dri/N1668_1_7  (
            .Z (_N10992_3),
            .I0 (_N10545),
            .I1 (_N10546),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I4 (_N10569),
            .ID (_N10568));
	// LUT = (I1&~I3&I4)|(I0&~I2&I4)|(I0&I1&I4)|(~I2&~I3)|(ID&I1&~I3) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1668_1_9  */ #(
            .INIT(32'b11111111010101011111111101010000))
        \u_touch_top/u_i2c_dri/N1668_1_9  (
            .Z (_N10992_1),
            .I0 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (_N10566),
            .I3 (_N10992_3),
            .I4 (_N11426_3));
	// LUT = (~I0&I4)|(I3)|(~I0&I2) ;

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N1668_4  */ #(
            .INIT(16'b1010100010101010))
        \u_touch_top/u_i2c_dri/N1668_4  (
            .Z (_N10344),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N10566));
	// LUT = (I0&~I3)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1668_5  */ #(
            .INIT(32'b10100000101010001010001010101010))
        \u_touch_top/u_i2c_dri/N1668_5  (
            .Z (_N10345),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [7] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N10568),
            .I4 (_N10569));
	// LUT = (I0&~I1&~I4)|(I0&I1&~I3)|(I0&I2) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1679_18_2  */ #(
            .INIT(32'b11111111111111101111111111111101))
        \u_touch_top/u_i2c_dri/N1679_18_2  (
            .Z (_N12029),
            .I0 (\u_touch_top/u_i2c_dri/N476 ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I4 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .ID (\u_touch_top/u_i2c_dri/cur_state_reg [1] ));
	// LUT = (~ID&~I4)|(I0&I4)|(I3)|(I2)|(I1) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1679_18_6  */ #(
            .INIT(32'b11111111111111111111111111111110))
        \u_touch_top/u_i2c_dri/N1679_18_6  (
            .Z (_N2517),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I4 (_N12029));
	// LUT = (I4)|(I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1679_22  */ #(
            .INIT(32'b00000000000001010000000000000001))
        \u_touch_top/u_i2c_dri/N1679_22  (
            .Z (_N2521),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I4 (\u_touch_top/u_i2c_dri/addr_t [0] ));
	// LUT = (~I0&~I2&~I3&I4)|(~I0&~I1&~I2&~I3) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1679_28_2  */ #(
            .INIT(32'b00000000001000100000000000110001))
        \u_touch_top/u_i2c_dri/N1679_28_2  (
            .Z (_N12037),
            .I0 (\u_touch_top/u_i2c_dri/data_wr_t [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I2 (\u_touch_top/u_i2c_dri/addr_t [1] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I4 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .ID (\u_touch_top/u_i2c_dri/cur_state_reg [3] ));
	// LUT = (~I1&I2&~I3&~I4)|(~ID&~I1&~I3&~I4)|(I0&~I1&~I3&I4) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1679_29  */ #(
            .INIT(32'b11010101100001011101000010000000))
        \u_touch_top/u_i2c_dri/N1679_29  (
            .Z (_N2528),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I1 (\u_touch_top/u_i2c_dri/addr_t [6] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N2521),
            .I4 (_N12037));
	// LUT = (~I0&~I2&I4)|(~I0&I2&I3)|(I0&I1&I2) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1679_44  */ #(
            .INIT(32'b11111111111110101111111111110010))
        \u_touch_top/u_i2c_dri/N1679_44  (
            .Z (_N2543),
            .I0 (_N2528),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .ID (_N11198_2));
	// LUT = (ID&~I1&~I4)|(I0&I4)|(I3)|(I2) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1679_53  */ #(
            .INIT(32'b10101010101010101111110100110001))
        \u_touch_top/u_i2c_dri/N1679_53  (
            .Z (_N2552),
            .I0 (\u_touch_top/slave_addr [4] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I2 (\u_touch_top/u_i2c_dri/addr_t [4] ),
            .I3 (\u_touch_top/u_i2c_dri/data_wr_t [1] ),
            .I4 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .ID (\u_touch_top/u_i2c_dri/cur_state_reg [3] ));
	// LUT = (I1&I3&~I4)|(~I1&I2&~I4)|(~ID&~I1&~I4)|(I0&I4) ;

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N1679_56  */ #(
            .INIT(4'b1101))
        \u_touch_top/u_i2c_dri/N1679_56  (
            .Z (_N2555),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I1 (\u_touch_top/u_i2c_dri/addr_t [5] ));
	// LUT = (I1)|(~I0) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1679_59  */ #(
            .INIT(32'b10101000101010111010100010101000))
        \u_touch_top/u_i2c_dri/N1679_59  (
            .Z (_N2558),
            .I0 (\u_touch_top/slave_addr [3] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I4 (_N2555));
	// LUT = (~I1&~I2&~I3&I4)|(I0&I2)|(I0&I1) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1679_61  */ #(
            .INIT(32'b00000000101110000000000010101010))
        \u_touch_top/u_i2c_dri/N1679_61  (
            .Z (_N2560),
            .I0 (\u_touch_top/slave_addr [4] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I2 (_N2552),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .ID (_N2558));
	// LUT = (ID&~I3&~I4)|(~I1&I2&~I3&I4)|(I0&I1&~I3&I4) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1679_69_2  */ #(
            .INIT(32'b00000000000001010000000000000001))
        \u_touch_top/u_i2c_dri/N1679_69_2  (
            .Z (_N12039),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I4 (\u_touch_top/u_i2c_dri/addr_t [6] ));
	// LUT = (~I0&~I2&~I3&I4)|(~I0&~I1&~I2&~I3) ;

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N1679_72  */ #(
            .INIT(16'b1100111111001101))
        \u_touch_top/u_i2c_dri/N1679_72  (
            .Z (_N2571),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I3 (\u_touch_top/u_i2c_dri/addr_t [7] ));
	// LUT = (~I2&I3)|(~I0&~I2)|(I1) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1679_75  */ #(
            .INIT(32'b00100010001000100000111000000010))
        \u_touch_top/u_i2c_dri/N1679_75  (
            .Z (_N2574),
            .I0 (_N12039),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [7] ),
            .I3 (\u_touch_top/u_i2c_dri/addr_t [6] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .ID (_N2571));
	// LUT = (I1&~I2&I3&~I4)|(ID&~I1&~I2&~I4)|(I0&~I1&I4) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1679_77  */ #(
            .INIT(32'b11101110111011101111011111000100))
        \u_touch_top/u_i2c_dri/N1679_77  (
            .Z (_N2576),
            .I0 (_N2560),
            .I1 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N2574),
            .I4 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .ID (\u_touch_top/u_i2c_dri/cur_state_reg [5] ));
	// LUT = (~I1&I3&~I4)|(I1&I4)|(I0&I4)|(I1&I2)|(~ID&I1) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1679_78  */ #(
            .INIT(32'b11111111111111011010101010101010))
        \u_touch_top/u_i2c_dri/N1679_78  (
            .Z (_N2577),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [1] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .ID (_N2576));
	// LUT = (ID&~I4)|(I3&I4)|(I2&I4)|(I1&I4)|(~I0&I4) ;

    GTP_MUX2LUT6 \u_touch_top/u_i2c_dri/N1679_79  (
            .Z (_N2578),
            .I0 (_N2577),
            .I1 (_N2543),
            .S (\u_touch_top/u_i2c_dri/cnt [4] ));

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N1679_101  */ #(
            .INIT(32'b10101011101010001010101110101000))
        \u_touch_top/u_i2c_dri/N1679_101  (
            .Z (_N11198_2),
            .I0 (\u_touch_top/bit_ctrl ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I3 (_N11198_5),
            .I4 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .ID (\u_touch_top/slave_addr [3] ));
	// LUT = (ID&I2&~I4)|(ID&I1&~I4)|(I0&I2&I4)|(I0&I1&I4)|(~I1&~I2&I3) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N1679_104  */ #(
            .INIT(32'b11110111110101011010001010000000))
        \u_touch_top/u_i2c_dri/N1679_104  (
            .Z (_N11198_5),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/data_wr_t [2] ),
            .I3 (\u_touch_top/u_i2c_dri/data_wr_t [3] ),
            .I4 (_N11198_6));
	// LUT = (~I0&I4)|(I0&~I1&I3)|(I0&I1&I2) ;

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N1679_105  */ #(
            .INIT(16'b1101110111110101))
        \u_touch_top/u_i2c_dri/N1679_105  (
            .Z (_N11198_6),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I1 (\u_touch_top/u_i2c_dri/addr_t [2] ),
            .I2 (\u_touch_top/u_i2c_dri/addr_t [3] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [2] ));
	// LUT = (I2&~I3)|(I1&I3)|(~I0) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N2079_1_2  */ #(
            .INIT(32'b00100010000000000010000000100000))
        \u_touch_top/u_i2c_dri/N2079_1_2  (
            .Z (_N12012),
            .I0 (_N10569),
            .I1 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .ID (_N10566));
	// LUT = (ID&~I1&I2&~I4)|(I0&~I1&I3&I4) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N2079_1_3  */ #(
            .INIT(32'b00000011000000100000000000000000))
        \u_touch_top/u_i2c_dri/N2079_1_3  (
            .Z (_N12013),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N10315),
            .I4 (_N10569));
	// LUT = (~I1&~I2&I3&I4)|(I0&~I1&~I2&I4) ;

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N2079_5_3  */ #(
            .INIT(16'b1111111111111110))
        \u_touch_top/u_i2c_dri/N2079_5_3  (
            .Z (_N10315),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [7] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N2079_28  */ #(
            .INIT(32'b11111111111111111111111111100000))
        \u_touch_top/u_i2c_dri/N2079_28  (
            .Z (\u_touch_top/u_i2c_dri/N1230 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I2 (\u_touch_top/u_i2c_dri/N1185 ),
            .I3 (\u_touch_top/u_i2c_dri/N1222 ),
            .I4 (_N10904_2));
	// LUT = (I4)|(I3)|(I1&I2)|(I0&I2) ;

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N2082_5  */ #(
            .INIT(16'b1111111000000000))
        \u_touch_top/u_i2c_dri/N2082_5  (
            .Z (_N10904_2),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I3 (\u_touch_top/u_i2c_dri/N1180 ));
	// LUT = (I2&I3)|(I1&I3)|(I0&I3) ;

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/N2434_6  */ #(
            .INIT(32'b11000000100000001000000010000000))
        \u_touch_top/u_i2c_dri/N2434_6  (
            .Z (\u_touch_top/u_i2c_dri/N2434 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (_N10566),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I4 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .ID (_N11792_3));
	// LUT = (ID&I1&I2&~I4)|(I1&I2&I3&I4)|(I0&I1&I2&I4) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N2868  */ #(
            .INIT(32'b10000000000000000000000000000000))
        \u_touch_top/u_i2c_dri/N2868_vname  (
            .Z (\u_touch_top/u_i2c_dri/N2868 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (_N10539),
            .I4 (_N10547));
    // defparam \u_touch_top/u_i2c_dri/N2868_vname .orig_name = \u_touch_top/u_i2c_dri/N2868 ;
	// LUT = I0&I1&I2&I3&I4 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N2917  */ #(
            .INIT(16'b0000100000000000))
        \u_touch_top/u_i2c_dri/N2917_vname  (
            .Z (\u_touch_top/u_i2c_dri/N2917 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N10566));
    // defparam \u_touch_top/u_i2c_dri/N2917_vname .orig_name = \u_touch_top/u_i2c_dri/N2917 ;
	// LUT = I0&I1&~I2&I3 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT2 /* \u_touch_top/u_i2c_dri/N2925  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_i2c_dri/N2925_vname  (
            .Z (\u_touch_top/u_i2c_dri/N2925 ),
            .I0 (\u_touch_top/i2c_exec ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [0] ));
    // defparam \u_touch_top/u_i2c_dri/N2925_vname .orig_name = \u_touch_top/u_i2c_dri/N2925 ;
	// LUT = I0&I1 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N3005  */ #(
            .INIT(32'b11001100110011101100110011001100))
        \u_touch_top/u_i2c_dri/N3005_vname  (
            .Z (\u_touch_top/u_i2c_dri/N3005 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I1 (\u_touch_top/u_i2c_dri/N2925 ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I3 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I4 (_N10569));
    // defparam \u_touch_top/u_i2c_dri/N3005_vname .orig_name = \u_touch_top/u_i2c_dri/N3005 ;
	// LUT = (I0&~I2&~I3&I4)|(I1) ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N3052  */ #(
            .INIT(16'b0000100000000000))
        \u_touch_top/u_i2c_dri/N3052_vname  (
            .Z (\u_touch_top/u_i2c_dri/N3052 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N10569));
    // defparam \u_touch_top/u_i2c_dri/N3052_vname .orig_name = \u_touch_top/u_i2c_dri/N3052 ;
	// LUT = I0&I1&~I2&I3 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/N3102  */ #(
            .INIT(16'b1000000000000000))
        \u_touch_top/u_i2c_dri/N3102_vname  (
            .Z (\u_touch_top/u_i2c_dri/N3102 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [2] ),
            .I3 (_N10569));
    // defparam \u_touch_top/u_i2c_dri/N3102_vname .orig_name = \u_touch_top/u_i2c_dri/N3102 ;
	// LUT = I0&I1&I2&I3 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N3152  */ #(
            .INIT(32'b00001000000000000000000000000000))
        \u_touch_top/u_i2c_dri/N3152_vname  (
            .Z (\u_touch_top/u_i2c_dri/N3152 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (_N10539),
            .I4 (_N10545));
    // defparam \u_touch_top/u_i2c_dri/N3152_vname .orig_name = \u_touch_top/u_i2c_dri/N3152 ;
	// LUT = I0&I1&~I2&I3&I4 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N3202  */ #(
            .INIT(32'b00001000000000000000000000000000))
        \u_touch_top/u_i2c_dri/N3202_vname  (
            .Z (\u_touch_top/u_i2c_dri/N3202 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (_N10539),
            .I4 (_N10547));
    // defparam \u_touch_top/u_i2c_dri/N3202_vname .orig_name = \u_touch_top/u_i2c_dri/N3202 ;
	// LUT = I0&I1&~I2&I3&I4 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N3252  */ #(
            .INIT(32'b00100000000000000000000000000000))
        \u_touch_top/u_i2c_dri/N3252_vname  (
            .Z (\u_touch_top/u_i2c_dri/N3252 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (_N10539),
            .I4 (_N10545));
    // defparam \u_touch_top/u_i2c_dri/N3252_vname .orig_name = \u_touch_top/u_i2c_dri/N3252 ;
	// LUT = I0&~I1&I2&I3&I4 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N3302  */ #(
            .INIT(32'b00100000000000000000000000000000))
        \u_touch_top/u_i2c_dri/N3302_vname  (
            .Z (\u_touch_top/u_i2c_dri/N3302 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (_N10539),
            .I4 (_N10547));
    // defparam \u_touch_top/u_i2c_dri/N3302_vname .orig_name = \u_touch_top/u_i2c_dri/N3302 ;
	// LUT = I0&~I1&I2&I3&I4 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/N3352  */ #(
            .INIT(32'b10000000000000000000000000000000))
        \u_touch_top/u_i2c_dri/N3352_vname  (
            .Z (\u_touch_top/u_i2c_dri/N3352 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cnt [4] ),
            .I3 (_N10539),
            .I4 (_N10545));
    // defparam \u_touch_top/u_i2c_dri/N3352_vname .orig_name = \u_touch_top/u_i2c_dri/N3352 ;
	// LUT = I0&I1&I2&I3&I4 ;
	// ../../rtl/touch/i2c_dri.v:227

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/ack  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/ack  (
            .Q (\u_touch_top/i2c_ack ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2434 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N3));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/addr_t[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/addr_t[0]  (
            .Q (\u_touch_top/u_i2c_dri/addr_t [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2925 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_addr [0] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/addr_t[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/addr_t[1]  (
            .Q (\u_touch_top/u_i2c_dri/addr_t [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2925 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_addr [1] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/addr_t[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/addr_t[2]  (
            .Q (\u_touch_top/u_i2c_dri/addr_t [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2925 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_addr [2] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/addr_t[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/addr_t[3]  (
            .Q (\u_touch_top/u_i2c_dri/addr_t [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2925 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_addr [3] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/addr_t[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/addr_t[4]  (
            .Q (\u_touch_top/u_i2c_dri/addr_t [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2925 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_addr [4] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/addr_t[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/addr_t[5]  (
            .Q (\u_touch_top/u_i2c_dri/addr_t [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2925 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_addr [5] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/addr_t[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/addr_t[6]  (
            .Q (\u_touch_top/u_i2c_dri/addr_t [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2925 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_addr [6] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/addr_t[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/addr_t[7]  (
            .Q (\u_touch_top/u_i2c_dri/addr_t [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2925 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_addr [7] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/clk_cnt[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/clk_cnt[0]  (
            .Q (\u_touch_top/u_i2c_dri/clk_cnt [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_sys_clk),
            .D (\u_touch_top/u_i2c_dri/clk_cnt[0]_inv ));
	// ../../rtl/touch/i2c_dri.v:86

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/clk_cnt[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/clk_cnt[1]  (
            .Q (\u_touch_top/u_i2c_dri/clk_cnt [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_sys_clk),
            .D (\u_touch_top/u_i2c_dri/N811 [1] ));
	// ../../rtl/touch/i2c_dri.v:86

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/clk_cnt[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/clk_cnt[2]  (
            .Q (\u_touch_top/u_i2c_dri/clk_cnt [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_sys_clk),
            .D (\u_touch_top/u_i2c_dri/N12 [2] ));
	// ../../rtl/touch/i2c_dri.v:86

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/clk_cnt[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/clk_cnt[3]  (
            .Q (\u_touch_top/u_i2c_dri/clk_cnt [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_sys_clk),
            .D (\u_touch_top/u_i2c_dri/N12 [3] ));
	// ../../rtl/touch/i2c_dri.v:86

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/clk_cnt[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/clk_cnt[4]  (
            .Q (\u_touch_top/u_i2c_dri/clk_cnt [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_sys_clk),
            .D (\u_touch_top/u_i2c_dri/N811 [4] ));
	// ../../rtl/touch/i2c_dri.v:86

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/clk_cnt[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/clk_cnt[5]  (
            .Q (\u_touch_top/u_i2c_dri/clk_cnt [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (nt_sys_clk),
            .D (\u_touch_top/u_i2c_dri/N811 [5] ));
	// ../../rtl/touch/i2c_dri.v:86

    GTP_LUT1 /* \u_touch_top/u_i2c_dri/clk_cnt[9:0]_inv  */ #(
            .INIT(2'b01))
        \u_touch_top/u_i2c_dri/clk_cnt[9:0]_inv  (
            .Z (\u_touch_top/u_i2c_dri/clk_cnt[0]_inv ),
            .I0 (\u_touch_top/u_i2c_dri/clk_cnt [0] ));
	// LUT = ~I0 ;

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cnt[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cnt[0]  (
            .Q (\u_touch_top/u_i2c_dri/cnt [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N552 [0] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cnt[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cnt[1]  (
            .Q (\u_touch_top/u_i2c_dri/cnt [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N552 [1] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cnt[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cnt[2]  (
            .Q (\u_touch_top/u_i2c_dri/cnt [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N552 [2] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cnt[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cnt[3]  (
            .Q (\u_touch_top/u_i2c_dri/cnt [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N552 [3] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cnt[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cnt[4]  (
            .Q (\u_touch_top/u_i2c_dri/cnt [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N552 [4] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cnt[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cnt[5]  (
            .Q (\u_touch_top/u_i2c_dri/cnt [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N552 [5] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cnt[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cnt[6]  (
            .Q (\u_touch_top/u_i2c_dri/cnt [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N552 [6] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_3  */ #(
            .INIT(16'b1111010001000100))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_3  (
            .Z (\u_touch_top/u_i2c_dri/_N2 ),
            .I0 (\u_touch_top/i2c_exec ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [7] ),
            .I3 (\u_touch_top/u_i2c_dri/st_done ));
	// LUT = (I2&I3)|(~I0&I1) ;
	// ../../rtl/touch/i2c_dri.v:110

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_6  */ #(
            .INIT(16'b1010000011101100))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_6  (
            .Z (\u_touch_top/u_i2c_dri/_N5 ),
            .I0 (\u_touch_top/i2c_exec ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [0] ),
            .I3 (\u_touch_top/u_i2c_dri/st_done ));
	// LUT = (I1&~I3)|(I0&I2) ;
	// ../../rtl/touch/i2c_dri.v:110

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_10  */ #(
            .INIT(32'b00100010000000001111000011110000))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_10  (
            .Z (\u_touch_top/u_i2c_dri/_N9 ),
            .I0 (\u_touch_top/bit_ctrl ),
            .I1 (\u_touch_top/i2c_ack ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I4 (\u_touch_top/u_i2c_dri/st_done ));
	// LUT = (I2&~I4)|(I0&~I1&I3&I4) ;
	// ../../rtl/touch/i2c_dri.v:110

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_16_3  */ #(
            .INIT(32'b00001111000001001010101010101010))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_16_3  (
            .Z (\u_touch_top/u_i2c_dri/_N15 ),
            .I0 (\u_touch_top/bit_ctrl ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I2 (\u_touch_top/i2c_ack ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I4 (\u_touch_top/u_i2c_dri/st_done ),
            .ID (\u_touch_top/u_i2c_dri/cur_state_reg [3] ));
	// LUT = (ID&~I4)|(~I2&I3&I4)|(~I0&I1&~I2&I4) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_20  */ #(
            .INIT(32'b00101010111111110010101000101010))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_20  (
            .Z (\u_touch_top/u_i2c_dri/_N19 ),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I1 (\u_touch_top/u_i2c_dri/reg_done ),
            .I2 (\u_touch_top/u_i2c_dri/st_done ),
            .I3 (\u_touch_top/u_i2c_dri/wr_flag ),
            .I4 (_N10558));
	// LUT = (~I3&I4)|(I0&~I2)|(I0&~I1) ;
	// ../../rtl/touch/i2c_dri.v:110

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_24  */ #(
            .INIT(32'b01000100111100000000000011110000))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_24  (
            .Z (\u_touch_top/u_i2c_dri/_N23 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I3 (\u_touch_top/u_i2c_dri/st_done ),
            .I4 (\u_touch_top/u_i2c_dri/wr_flag ));
	// LUT = (~I0&I1&I3&I4)|(I2&~I3) ;
	// ../../rtl/touch/i2c_dri.v:110

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_28  */ #(
            .INIT(32'b01010000110111001100110011001100))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_28  (
            .Z (\u_touch_top/u_i2c_dri/_N27 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .I3 (\u_touch_top/u_i2c_dri/reg_done ),
            .I4 (\u_touch_top/u_i2c_dri/st_done ));
	// LUT = (I1&~I4)|(~I0&I2&I4)|(I1&~I3) ;
	// ../../rtl/touch/i2c_dri.v:110

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_59_3  */ #(
            .INIT(32'b11101110111010101010101010101010))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_59_3  (
            .Z (\u_touch_top/u_i2c_dri/_N39 ),
            .I0 (_N12002),
            .I1 (\u_touch_top/u_i2c_dri/reg_done ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .I4 (\u_touch_top/u_i2c_dri/st_done ),
            .ID (\u_touch_top/u_i2c_dri/cur_state_reg [7] ));
	// LUT = (ID&~I4)|(I1&I3&I4)|(I1&I2&I4)|(I0&I4) ;

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_61_2  */ #(
            .INIT(32'b10101010101010101010101010101000))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_61_2  (
            .Z (_N12002),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .I3 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I4 (\u_touch_top/u_i2c_dri/cur_state_reg [5] ));
	// LUT = (I0&I4)|(I0&I3)|(I0&I2)|(I0&I1) ;

    GTP_LUT3 /* \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_70  */ #(
            .INIT(8'b00001000))
        \u_touch_top/u_i2c_dri/cur_state_fsm[7:0]_70  (
            .Z (_N10532),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ));
	// LUT = I0&I1&~I2 ;

(* syn_encoding="onehot" *)    GTP_DFF_P /* \u_touch_top/u_i2c_dri/cur_state_reg[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b1))
        \u_touch_top/u_i2c_dri/cur_state_reg[0]  (
            .Q (\u_touch_top/u_i2c_dri/cur_state_reg [0] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/_N2 ),
            .P (\u_lcd_rgb_char/u_binary2bcd_x/N0 ));
	// ../../rtl/touch/i2c_dri.v:110

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cur_state_reg[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cur_state_reg[1]  (
            .Q (\u_touch_top/u_i2c_dri/cur_state_reg [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/_N5 ));
	// ../../rtl/touch/i2c_dri.v:110

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cur_state_reg[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cur_state_reg[2]  (
            .Q (\u_touch_top/u_i2c_dri/cur_state_reg [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/_N9 ));
	// ../../rtl/touch/i2c_dri.v:110

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cur_state_reg[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cur_state_reg[3]  (
            .Q (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/_N15 ));
	// ../../rtl/touch/i2c_dri.v:110

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cur_state_reg[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cur_state_reg[4]  (
            .Q (\u_touch_top/u_i2c_dri/cur_state_reg [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/_N19 ));
	// ../../rtl/touch/i2c_dri.v:110

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cur_state_reg[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cur_state_reg[5]  (
            .Q (\u_touch_top/u_i2c_dri/cur_state_reg [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/_N23 ));
	// ../../rtl/touch/i2c_dri.v:110

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cur_state_reg[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cur_state_reg[6]  (
            .Q (\u_touch_top/u_i2c_dri/cur_state_reg [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/_N27 ));
	// ../../rtl/touch/i2c_dri.v:110

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_i2c_dri/cur_state_reg[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/cur_state_reg[7]  (
            .Q (\u_touch_top/u_i2c_dri/cur_state_reg [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/_N39 ));
	// ../../rtl/touch/i2c_dri.v:110

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_r[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_r[0]  (
            .Q (\u_touch_top/u_i2c_dri/data_r [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2868 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N3));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_r[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_r[1]  (
            .Q (\u_touch_top/u_i2c_dri/data_r [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3352 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N3));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_r[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_r[2]  (
            .Q (\u_touch_top/u_i2c_dri/data_r [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3302 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N3));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_r[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_r[3]  (
            .Q (\u_touch_top/u_i2c_dri/data_r [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3252 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N3));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_r[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_r[4]  (
            .Q (\u_touch_top/u_i2c_dri/data_r [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3202 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N3));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_r[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_r[5]  (
            .Q (\u_touch_top/u_i2c_dri/data_r [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3152 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N3));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_r[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_r[6]  (
            .Q (\u_touch_top/u_i2c_dri/data_r [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3102 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N3));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_r[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_r[7]  (
            .Q (\u_touch_top/u_i2c_dri/data_r [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3052 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N3));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_wr_t[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_wr_t[1]  (
            .Q (\u_touch_top/u_i2c_dri/data_wr_t [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3005 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_w [1] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_wr_t[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_wr_t[2]  (
            .Q (\u_touch_top/u_i2c_dri/data_wr_t [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3005 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_w [2] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/data_wr_t[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/data_wr_t[3]  (
            .Q (\u_touch_top/u_i2c_dri/data_wr_t [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N3005 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_w [3] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_PE /* \u_touch_top/u_i2c_dri/dri_clk  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b1))
        \u_touch_top/u_i2c_dri/dri_clk  (
            .Q (\u_touch_top/dri_clk ),
            .CE (1'b1),
            .CLK (nt_sys_clk),
            .D (_N11806),
            .P (\u_lcd_rgb_char/u_binary2bcd_x/N0 ));
	// ../../rtl/touch/i2c_dri.v:86

    GTP_LUT4 /* \u_touch_top/u_i2c_dri/dri_clk_ce_mux  */ #(
            .INIT(16'b0110101010101010))
        \u_touch_top/u_i2c_dri/dri_clk_ce_mux  (
            .Z (_N11806),
            .I0 (\u_touch_top/dri_clk ),
            .I1 (\u_touch_top/u_i2c_dri/clk_cnt [0] ),
            .I2 (\u_touch_top/u_i2c_dri/clk_cnt [5] ),
            .I3 (_N12050));
	// LUT = (I0&~I3)|(~I0&I1&I2&I3)|(I0&~I2)|(I0&~I1) ;

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/i2c_data_r[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/i2c_data_r[0]  (
            .Q (\u_touch_top/i2c_data_r [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2917 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/data_r [0] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/i2c_data_r[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/i2c_data_r[1]  (
            .Q (\u_touch_top/i2c_data_r [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2917 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/data_r [1] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/i2c_data_r[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/i2c_data_r[2]  (
            .Q (\u_touch_top/i2c_data_r [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2917 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/data_r [2] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/i2c_data_r[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/i2c_data_r[3]  (
            .Q (\u_touch_top/i2c_data_r [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2917 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/data_r [3] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/i2c_data_r[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/i2c_data_r[4]  (
            .Q (\u_touch_top/i2c_data_r [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2917 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/data_r [4] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/i2c_data_r[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/i2c_data_r[5]  (
            .Q (\u_touch_top/i2c_data_r [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2917 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/data_r [5] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/i2c_data_r[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/i2c_data_r[6]  (
            .Q (\u_touch_top/i2c_data_r [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2917 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/data_r [6] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/i2c_data_r[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/i2c_data_r[7]  (
            .Q (\u_touch_top/i2c_data_r [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2917 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/data_r [7] ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/i2c_done  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/i2c_done  (
            .Q (\u_touch_top/i2c_done ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (1'b1),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N11814));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/i2c_done_ce_mux  */ #(
            .INIT(32'b00110010001000100010001000100010))
        \u_touch_top/u_i2c_dri/i2c_done_ce_mux  (
            .Z (_N11814),
            .I0 (\u_touch_top/i2c_done ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [0] ),
            .I2 (\u_touch_top/u_i2c_dri/cur_state_reg [7] ),
            .I3 (_N10548),
            .I4 (_N10568));
	// LUT = (~I1&I2&I3&I4)|(I0&~I1) ;

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/once_byte_done  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/once_byte_done  (
            .Q (\u_touch_top/once_byte_done ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N558 ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/reg_cnt[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/reg_cnt[0]  (
            .Q (\u_touch_top/u_i2c_dri/reg_cnt [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N814 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N815 [0] ));
	// ../../rtl/touch/i2c_dri.v:100

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/reg_cnt[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/reg_cnt[1]  (
            .Q (\u_touch_top/u_i2c_dri/reg_cnt [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N814 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N815 [1] ));
	// ../../rtl/touch/i2c_dri.v:100

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/reg_cnt[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/reg_cnt[2]  (
            .Q (\u_touch_top/u_i2c_dri/reg_cnt [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N814 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N815 [2] ));
	// ../../rtl/touch/i2c_dri.v:100

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/reg_cnt[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/reg_cnt[3]  (
            .Q (\u_touch_top/u_i2c_dri/reg_cnt [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N814 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N815 [3] ));
	// ../../rtl/touch/i2c_dri.v:100

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/reg_cnt[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/reg_cnt[4]  (
            .Q (\u_touch_top/u_i2c_dri/reg_cnt [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N814 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N815 [4] ));
	// ../../rtl/touch/i2c_dri.v:100

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/reg_cnt[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/reg_cnt[5]  (
            .Q (\u_touch_top/u_i2c_dri/reg_cnt [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N814 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N815 [5] ));
	// ../../rtl/touch/i2c_dri.v:100

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/reg_cnt[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/reg_cnt[6]  (
            .Q (\u_touch_top/u_i2c_dri/reg_cnt [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N814 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N815 [6] ));
	// ../../rtl/touch/i2c_dri.v:100

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/reg_cnt[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/reg_cnt[7]  (
            .Q (\u_touch_top/u_i2c_dri/reg_cnt [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N814 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N815 [7] ));
	// ../../rtl/touch/i2c_dri.v:100

    GTP_DFF_PE /* \u_touch_top/u_i2c_dri/scl  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b1))
        \u_touch_top/u_i2c_dri/scl  (
            .Q (nt_touch_scl),
            .CE (\u_touch_top/u_i2c_dri/N1227 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N1232 ),
            .P (\u_lcd_rgb_char/u_binary2bcd_x/N0 ));
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_PE /* \u_touch_top/u_i2c_dri/sda_dir  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b1))
        \u_touch_top/u_i2c_dri/sda_dir_vname  (
            .Q (\u_touch_top/u_i2c_dri/sda_dir ),
            .CE (1'b1),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N11813),
            .P (\u_lcd_rgb_char/u_binary2bcd_x/N0 ));
    // defparam \u_touch_top/u_i2c_dri/sda_dir_vname .orig_name = \u_touch_top/u_i2c_dri/sda_dir ;
	// ../../rtl/touch/i2c_dri.v:206

    GTP_LUT5 /* \u_touch_top/u_i2c_dri/sda_dir_ce_mux  */ #(
            .INIT(32'b00110011001100110011001100110010))
        \u_touch_top/u_i2c_dri/sda_dir_ce_mux  (
            .Z (_N11813),
            .I0 (\u_touch_top/u_i2c_dri/cur_state_reg [0] ),
            .I1 (\u_touch_top/u_i2c_dri/N2082 ),
            .I2 (\u_touch_top/u_i2c_dri/sda_dir ),
            .I3 (_N12012),
            .I4 (_N12013));
	// LUT = (~I1&I4)|(~I1&I3)|(~I1&I2)|(I0&~I1) ;

    GTP_LUT1 /* \u_touch_top/u_i2c_dri/sda_dir_inv  */ #(
            .INIT(2'b01))
        \u_touch_top/u_i2c_dri/sda_dir_inv_vname  (
            .Z (\u_touch_top/u_i2c_dri/sda_dir_inv ),
            .I0 (\u_touch_top/u_i2c_dri/sda_dir ));
    // defparam \u_touch_top/u_i2c_dri/sda_dir_inv_vname .orig_name = \u_touch_top/u_i2c_dri/sda_dir_inv ;
	// LUT = ~I0 ;

    GTP_DFF_PE /* \u_touch_top/u_i2c_dri/sda_out  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b1))
        \u_touch_top/u_i2c_dri/sda_out_vname  (
            .Q (\u_touch_top/u_i2c_dri/sda_out ),
            .CE (1'b1),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N11812),
            .P (\u_lcd_rgb_char/u_binary2bcd_x/N0 ));
    // defparam \u_touch_top/u_i2c_dri/sda_out_vname .orig_name = \u_touch_top/u_i2c_dri/sda_out ;
	// ../../rtl/touch/i2c_dri.v:206

    GTP_LUT5M /* \u_touch_top/u_i2c_dri/sda_out_ce_mux  */ #(
            .INIT(32'b10101010101010101111110111101100))
        \u_touch_top/u_i2c_dri/sda_out_ce_mux  (
            .Z (_N11812),
            .I0 (\u_touch_top/u_i2c_dri/sda_out ),
            .I1 (\u_touch_top/u_i2c_dri/cnt [6] ),
            .I2 (_N2517),
            .I3 (_N2578),
            .I4 (\u_touch_top/u_i2c_dri/N1668 ),
            .ID (\u_touch_top/u_i2c_dri/cnt [5] ));
	// LUT = (~ID&I3&~I4)|(ID&I2&~I4)|(I1&~I4)|(I0&I4) ;

    GTP_DFF_C /* \u_touch_top/u_i2c_dri/st_done  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/st_done_vname  (
            .Q (\u_touch_top/u_i2c_dri/st_done ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_i2c_dri/N557 ));
    // defparam \u_touch_top/u_i2c_dri/st_done_vname .orig_name = \u_touch_top/u_i2c_dri/st_done ;
	// ../../rtl/touch/i2c_dri.v:206

    GTP_DFF_CE /* \u_touch_top/u_i2c_dri/wr_flag  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_i2c_dri/wr_flag_vname  (
            .Q (\u_touch_top/u_i2c_dri/wr_flag ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_i2c_dri/N2925 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_rh_wl ));
    // defparam \u_touch_top/u_i2c_dri/wr_flag_vname .orig_name = \u_touch_top/u_i2c_dri/wr_flag ;
	// ../../rtl/touch/i2c_dri.v:206

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_0  */ #(
            .INIT(32'b11001100110011000000000000000000), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("FALSE"), 
            .I4_TO_CARRY("FALSE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_0  (
            .COUT (_N655),
            .Z (),
            .CIN (),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [0] ),
            .I2 (),
            .I3 (),
            .I4 (),
            .ID ());
	// LUT = I1 ;
	// CARRY = (1'b0) ? CIN : (I1) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_1  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_1  (
            .COUT (_N656),
            .Z (\u_touch_top/u_touch_dri/N559 [1] ),
            .CIN (_N655),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [1] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_2  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_2  (
            .COUT (_N657),
            .Z (\u_touch_top/u_touch_dri/N559 [2] ),
            .CIN (_N656),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [2] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_3  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_3  (
            .COUT (_N658),
            .Z (\u_touch_top/u_touch_dri/N559 [3] ),
            .CIN (_N657),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [3] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_4  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_4  (
            .COUT (_N659),
            .Z (\u_touch_top/u_touch_dri/N559 [4] ),
            .CIN (_N658),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [4] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_5  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_5  (
            .COUT (_N660),
            .Z (\u_touch_top/u_touch_dri/N559 [5] ),
            .CIN (_N659),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [5] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_6  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_6  (
            .COUT (_N661),
            .Z (\u_touch_top/u_touch_dri/N559 [6] ),
            .CIN (_N660),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [6] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_7  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_7  (
            .COUT (_N662),
            .Z (\u_touch_top/u_touch_dri/N559 [7] ),
            .CIN (_N661),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [7] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_8  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_8  (
            .COUT (_N663),
            .Z (\u_touch_top/u_touch_dri/N559 [8] ),
            .CIN (_N662),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [8] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_9  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_9  (
            .COUT (_N664),
            .Z (\u_touch_top/u_touch_dri/N559 [9] ),
            .CIN (_N663),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [9] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_10  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_10  (
            .COUT (_N665),
            .Z (\u_touch_top/u_touch_dri/N559 [10] ),
            .CIN (_N664),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [10] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_11  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_11  (
            .COUT (_N666),
            .Z (\u_touch_top/u_touch_dri/N559 [11] ),
            .CIN (_N665),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [11] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_12  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_12  (
            .COUT (_N667),
            .Z (\u_touch_top/u_touch_dri/N559 [12] ),
            .CIN (_N666),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [12] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_13  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_13  (
            .COUT (_N668),
            .Z (\u_touch_top/u_touch_dri/N559 [13] ),
            .CIN (_N667),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [13] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_14  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_14  (
            .COUT (_N669),
            .Z (\u_touch_top/u_touch_dri/N559 [14] ),
            .CIN (_N668),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [14] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_15  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_15  (
            .COUT (_N670),
            .Z (\u_touch_top/u_touch_dri/N559 [15] ),
            .CIN (_N669),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [15] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_16  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_16  (
            .COUT (_N671),
            .Z (\u_touch_top/u_touch_dri/N559 [16] ),
            .CIN (_N670),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [16] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_17  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_17  (
            .COUT (_N672),
            .Z (\u_touch_top/u_touch_dri/N559 [17] ),
            .CIN (_N671),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [17] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_18  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_18  (
            .COUT (_N673),
            .Z (\u_touch_top/u_touch_dri/N559 [18] ),
            .CIN (_N672),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [18] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5CARRY /* \u_touch_top/u_touch_dri/N4_1_19  */ #(
            .INIT(32'b01100000011000001100110011001100), 
            .ID_TO_LUT("FALSE"), 
            .CIN_TO_LUT("TRUE"), 
            .I4_TO_CARRY("TRUE"), 
            .I4_TO_LUT("FALSE"))
        \u_touch_top/u_touch_dri/N4_1_19  (
            .COUT (),
            .Z (\u_touch_top/u_touch_dri/N559 [19] ),
            .CIN (_N673),
            .I0 (),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [19] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I3 (),
            .I4 (1'b0),
            .ID ());
	// LUT = (CIN&~I1&I2)|(~CIN&I1&I2) ;
	// CARRY = (I1) ? CIN : (I4) ;
	// ../../rtl/touch/touch_dri.v:107

    GTP_LUT5M /* \u_touch_top/u_touch_dri/N54_8[2]  */ #(
            .INIT(32'b01010101000000001111000100001100))
        \u_touch_top/u_touch_dri/N54_8[2]  (
            .Z (_N4964),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [4] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [3] ),
            .I3 (\u_touch_top/u_touch_dri/st_done ),
            .I4 (\u_touch_top/u_touch_dri/cur_state_reg [2] ),
            .ID (\u_touch_top/u_touch_dri/cur_state_reg [5] ));
	// LUT = (I1&~I2&~I3&~I4)|(I2&I3&~I4)|(~ID&~I1&I3&~I4)|(~I0&I3&I4) ;

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N54_8[3]_1  */ #(
            .INIT(4'b0001))
        \u_touch_top/u_touch_dri/N54_8[3]_1  (
            .Z (_N10511),
            .I0 (\u_touch_top/u_touch_dri/cur_state_reg [3] ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [2] ));
	// LUT = ~I0&~I1 ;

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N54_10[1]  */ #(
            .INIT(8'b10100100))
        \u_touch_top/u_touch_dri/N54_10[1]  (
            .Z (\u_touch_top/u_touch_dri/next_state [1] ),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
	// LUT = (~I0&I1&~I2)|(I0&I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N54_10[2]  */ #(
            .INIT(16'b0000000010100100))
        \u_touch_top/u_touch_dri/N54_10[2]  (
            .Z (\u_touch_top/u_touch_dri/next_state [2] ),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [2] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I3 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
	// LUT = (~I0&I1&~I2&~I3)|(I0&I2&~I3) ;

    GTP_LUT5M /* \u_touch_top/u_touch_dri/N54_10[3]_2  */ #(
            .INIT(32'b00000000000010000000000000000010))
        \u_touch_top/u_touch_dri/N54_10[3]_2  (
            .Z (\u_touch_top/u_touch_dri/next_state [3] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [2] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I3 (\u_touch_top/u_touch_dri/cur_state_reg [0] ),
            .I4 (\u_touch_top/u_touch_dri/st_done ),
            .ID (\u_touch_top/u_touch_dri/cur_state_reg [3] ));
	// LUT = (ID&~I1&~I2&~I3&~I4)|(I0&I1&~I2&~I3&I4) ;

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N54_10[4]_2  */ #(
            .INIT(8'b00010000))
        \u_touch_top/u_touch_dri/N54_10[4]_2  (
            .Z (\u_touch_top/u_touch_dri/next_state [4] ),
            .I0 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [0] ),
            .I2 (_N4964));
	// LUT = ~I0&~I1&I2 ;

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N54_10[5]_2  */ #(
            .INIT(4'b0001))
        \u_touch_top/u_touch_dri/N54_10[5]_2  (
            .Z (_N11987),
            .I0 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
	// LUT = ~I0&~I1 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N54_10[5]_3  */ #(
            .INIT(32'b10100100000000000000000000000000))
        \u_touch_top/u_touch_dri/N54_10[5]_3  (
            .Z (\u_touch_top/u_touch_dri/next_state [5] ),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [5] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [4] ),
            .I3 (_N10511),
            .I4 (_N11987));
	// LUT = (~I0&I1&~I2&I3&I4)|(I0&I2&I3&I4) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N54_10[6]_4  */ #(
            .INIT(32'b00001001000000000000000000000000))
        \u_touch_top/u_touch_dri/N54_10[6]_4  (
            .Z (\u_touch_top/u_touch_dri/next_state [6] ),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [5] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [4] ),
            .I3 (_N10511),
            .I4 (_N11987));
	// LUT = (~I0&~I1&~I2&I3&I4)|(I0&I1&~I2&I3&I4) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N70_mux18_2  */ #(
            .INIT(16'b0000000000011111))
        \u_touch_top/u_touch_dri/N70_mux18_2  (
            .Z (_N11972),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [1] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [2] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [3] ),
            .I3 (\u_touch_top/u_touch_dri/cnt_time [9] ));
	// LUT = (~I2&~I3)|(~I0&~I1&~I3) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N70_mux18_6  */ #(
            .INIT(32'b00010000000000000000000000000000))
        \u_touch_top/u_touch_dri/N70_mux18_6  (
            .Z (\u_touch_top/u_touch_dri/N70 ),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [10] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [13] ),
            .I2 (_N10520),
            .I3 (_N10560),
            .I4 (_N11972));
	// LUT = ~I0&~I1&I2&I3&I4 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N78_mux6_2  */ #(
            .INIT(32'b00000000000000011111111111111111))
        \u_touch_top/u_touch_dri/N78_mux6_2  (
            .Z (_N12192),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [4] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [5] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [6] ),
            .I3 (\u_touch_top/u_touch_dri/cnt_time [7] ),
            .I4 (\u_touch_top/u_touch_dri/cnt_time [9] ));
	// LUT = (~I4)|(~I0&~I1&~I2&~I3) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N78_mux8  */ #(
            .INIT(32'b00000000000011110000000000000111))
        \u_touch_top/u_touch_dri/N78_mux8  (
            .Z (_N574),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [8] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [10] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [11] ),
            .I3 (\u_touch_top/u_touch_dri/cnt_time [12] ),
            .I4 (_N12192));
	// LUT = (~I2&~I3&I4)|(~I1&~I2&~I3)|(~I0&~I2&~I3) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N78_mux8_4  */ #(
            .INIT(16'b0000000000000001))
        \u_touch_top/u_touch_dri/N78_mux8_4  (
            .Z (_N10457),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [16] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [17] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [18] ),
            .I3 (\u_touch_top/u_touch_dri/cnt_time [19] ));
	// LUT = ~I0&~I1&~I2&~I3 ;

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N113  */ #(
            .INIT(4'b1110))
        \u_touch_top/u_touch_dri/N113  (
            .Z (\u_touch_top/u_touch_dri/N1629 [9] ),
            .I0 (\u_lcd_rgb_char/u_clk_div/N40 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N152_26  */ #(
            .INIT(16'b1000000000000111))
        \u_touch_top/u_touch_dri/N152_26  (
            .Z (_N10246),
            .I0 (\u_touch_top/u_touch_dri/chip_version [0] ),
            .I1 (\u_touch_top/u_touch_dri/chip_version [1] ),
            .I2 (\u_touch_top/u_touch_dri/chip_version [12] ),
            .I3 (\u_touch_top/u_touch_dri/chip_version [13] ));
	// LUT = (~I1&~I2&~I3)|(~I0&~I2&~I3)|(I0&I1&I2&I3) ;

    GTP_LUT1 /* \u_touch_top/u_touch_dri/N166_1  */ #(
            .INIT(2'b01))
        \u_touch_top/u_touch_dri/N166_1  (
            .Z (\u_touch_top/u_touch_dri/N166 ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ));
	// LUT = ~I0 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N296  */ #(
            .INIT(32'b00000000001111100000000000000000))
        \u_touch_top/u_touch_dri/N296_vname  (
            .Z (\u_touch_top/u_touch_dri/N296 ),
            .I0 (\u_touch_top/i2c_data_r [0] ),
            .I1 (\u_touch_top/i2c_data_r [1] ),
            .I2 (\u_touch_top/i2c_data_r [2] ),
            .I3 (\u_touch_top/i2c_data_r [3] ),
            .I4 (_N10844));
    // defparam \u_touch_top/u_touch_dri/N296_vname .orig_name = \u_touch_top/u_touch_dri/N296 ;
	// LUT = (I1&~I2&~I3&I4)|(~I1&I2&~I3&I4)|(I0&~I1&~I3&I4) ;

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N296_1  */ #(
            .INIT(4'b1110))
        \u_touch_top/u_touch_dri/N296_1  (
            .Z (_N10844),
            .I0 (\u_touch_top/i2c_data_r [7] ),
            .I1 (\u_touch_top/u_touch_dri/ft_flag ));
	// LUT = (I1)|(I0) ;

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[0]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[0]  (
            .Z (\u_touch_top/u_touch_dri/N376 [0] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [0] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [8] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[1]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[1]  (
            .Z (\u_touch_top/u_touch_dri/N376 [1] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [1] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [9] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[2]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[2]  (
            .Z (\u_touch_top/u_touch_dri/N376 [2] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [2] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [10] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[3]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[3]  (
            .Z (\u_touch_top/u_touch_dri/N376 [3] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [3] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [11] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[4]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[4]  (
            .Z (\u_touch_top/u_touch_dri/N376 [4] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [4] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [12] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[5]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[5]  (
            .Z (\u_touch_top/u_touch_dri/N376 [5] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [5] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [13] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[6]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[6]  (
            .Z (\u_touch_top/u_touch_dri/N376 [6] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [6] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [14] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[7]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[7]  (
            .Z (\u_touch_top/u_touch_dri/N376 [7] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [7] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [15] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[8]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[8]  (
            .Z (\u_touch_top/u_touch_dri/N376 [8] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [8] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [0] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[9]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[9]  (
            .Z (\u_touch_top/u_touch_dri/N376 [9] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [9] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [1] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[10]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[10]  (
            .Z (\u_touch_top/u_touch_dri/N376 [10] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [10] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [2] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N376[11]  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/N376[11]  (
            .Z (\u_touch_top/u_touch_dri/N376 [11] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [11] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [3] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N376[12]_1  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/N376[12]_1  (
            .Z (\u_touch_top/u_touch_dri/N376 [12] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [12] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N376[13]_1  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/N376[13]_1  (
            .Z (\u_touch_top/u_touch_dri/N376 [13] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [13] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N376[14]_1  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/N376[14]_1  (
            .Z (\u_touch_top/u_touch_dri/N376 [14] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [14] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N376[15]_1  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/N376[15]_1  (
            .Z (\u_touch_top/u_touch_dri/N376 [15] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [15] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[0]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[0]  (
            .Z (\u_touch_top/u_touch_dri/N377 [0] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [8] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [0] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[1]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[1]  (
            .Z (\u_touch_top/u_touch_dri/N377 [1] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [9] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [1] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[2]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[2]  (
            .Z (\u_touch_top/u_touch_dri/N377 [2] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [10] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [2] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[3]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[3]  (
            .Z (\u_touch_top/u_touch_dri/N377 [3] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [11] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [3] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[4]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[4]  (
            .Z (\u_touch_top/u_touch_dri/N377 [4] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [12] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [4] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[5]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[5]  (
            .Z (\u_touch_top/u_touch_dri/N377 [5] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [13] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [5] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[6]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[6]  (
            .Z (\u_touch_top/u_touch_dri/N377 [6] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [14] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [6] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[7]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[7]  (
            .Z (\u_touch_top/u_touch_dri/N377 [7] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [15] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [7] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[8]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[8]  (
            .Z (\u_touch_top/u_touch_dri/N377 [8] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [0] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [8] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[9]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[9]  (
            .Z (\u_touch_top/u_touch_dri/N377 [9] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [1] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [9] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[10]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[10]  (
            .Z (\u_touch_top/u_touch_dri/N377 [10] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [2] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [10] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N377[11]  */ #(
            .INIT(8'b11011000))
        \u_touch_top/u_touch_dri/N377[11]  (
            .Z (\u_touch_top/u_touch_dri/N377 [11] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_x_coord_t [3] ),
            .I2 (\u_touch_top/u_touch_dri/tp_y_coord_t [11] ));
	// LUT = (~I0&I2)|(I0&I1) ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N377[12]_1  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/N377[12]_1  (
            .Z (\u_touch_top/u_touch_dri/N377 [12] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_y_coord_t [12] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N377[13]_1  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/N377[13]_1  (
            .Z (\u_touch_top/u_touch_dri/N377 [13] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_y_coord_t [13] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N377[14]_1  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/N377[14]_1  (
            .Z (\u_touch_top/u_touch_dri/N377 [14] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_y_coord_t [14] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N377[15]_1  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/N377[15]_1  (
            .Z (\u_touch_top/u_touch_dri/N377 [15] ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/tp_y_coord_t [15] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/touch/touch_dri.v:483

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N390_18_2  */ #(
            .INIT(32'b00000000000000000000000000000100))
        \u_touch_top/u_touch_dri/N390_18_2  (
            .Z (_N11979),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [5] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [6] ));
	// LUT = ~I0&I1&~I2&~I3&~I4 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N390_20_4  */ #(
            .INIT(32'b00000000000010000000000000000000))
        \u_touch_top/u_touch_dri/N390_20_4  (
            .Z (_N5000),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I1 (\u_touch_top/u_touch_dri/touch_valid ),
            .I2 (\u_touch_top/u_touch_dri/next_state [5] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [6] ),
            .I4 (_N10441));
	// LUT = I0&I1&~I2&~I3&I4 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N390_23  */ #(
            .INIT(32'b00000000111111110000001000000000))
        \u_touch_top/u_touch_dri/N390_23  (
            .Z (_N5003),
            .I0 (\u_touch_top/once_byte_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I2 (\u_touch_top/u_touch_dri/N1610 ),
            .I3 (\u_touch_top/u_touch_dri/next_state [5] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [6] ));
	// LUT = (I0&~I1&~I2&I3&~I4)|(~I3&I4) ;

    GTP_LUT5M /* \u_touch_top/u_touch_dri/N390_25  */ #(
            .INIT(32'b10101010000000001011100010111000))
        \u_touch_top/u_touch_dri/N390_25  (
            .Z (_N5005),
            .I0 (_N11979),
            .I1 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I2 (_N5003),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [7] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [3] ),
            .ID (_N5000));
	// LUT = (~I1&I2&~I4)|(ID&I1&~I4)|(I0&I3&I4) ;

    GTP_LUT5M /* \u_touch_top/u_touch_dri/N390_27  */ #(
            .INIT(32'b00100010000000001110001000100010))
        \u_touch_top/u_touch_dri/N390_27  (
            .Z (_N5007),
            .I0 (\u_touch_top/u_touch_dri/N474 ),
            .I1 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I3 (_N10521),
            .I4 (\u_touch_top/u_touch_dri/next_state [1] ),
            .ID (_N5005));
	// LUT = (I1&I2&I3&~I4)|(ID&~I1&~I4)|(I0&~I1&I3&I4) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N390_28  */ #(
            .INIT(16'b1101111100010000))
        \u_touch_top/u_touch_dri/N390_28  (
            .Z (\u_touch_top/u_touch_dri/N390 ),
            .I0 (\u_touch_top/u_touch_dri/N70 ),
            .I1 (\u_touch_top/u_touch_dri/st_done ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [0] ),
            .I3 (_N5007));
	// LUT = (~I2&I3)|(I1&I3)|(~I0&~I1&I2) ;

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N390_30  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/N390_30  (
            .Z (_N10441),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ));
	// LUT = ~I0&I1 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N390_73  */ #(
            .INIT(32'b00000000000001000000000000000000))
        \u_touch_top/u_touch_dri/N390_73  (
            .Z (_N11890),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [4] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [5] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [8] ),
            .I3 (\u_touch_top/u_touch_dri/cnt_time [12] ),
            .I4 (_N10517));
	// LUT = ~I0&I1&~I2&~I3&I4 ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N394_1_and[0][1]  */ #(
            .INIT(16'b0000000001000000))
        \u_touch_top/u_touch_dri/N394_1_and[0][1]  (
            .Z (_N9388),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [7] ));
	// LUT = ~I0&I1&I2&~I3 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N394_1_or[0]_7  */ #(
            .INIT(32'b11111111111111111110111111101110))
        \u_touch_top/u_touch_dri/N394_1_or[0]_7  (
            .Z (\u_touch_top/u_touch_dri/N394 ),
            .I0 (\u_touch_top/u_touch_dri/N945 ),
            .I1 (\u_touch_top/u_touch_dri/N1206 ),
            .I2 (\u_touch_top/u_touch_dri/N1610 ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I4 (_N9388));
	// LUT = (I4)|(~I2&I3)|(I1)|(I0) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N474_5  */ #(
            .INIT(32'b10000000000000000000000000000000))
        \u_touch_top/u_touch_dri/N474_5  (
            .Z (_N11935),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [11] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [14] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [15] ),
            .I3 (_N10457),
            .I4 (_N11890));
	// LUT = I0&I1&I2&I3&I4 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N474_7  */ #(
            .INIT(32'b00000010000000000000000000000000))
        \u_touch_top/u_touch_dri/N474_7  (
            .Z (\u_touch_top/u_touch_dri/N474 ),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [6] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [7] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [10] ),
            .I3 (\u_touch_top/u_touch_dri/cnt_time [13] ),
            .I4 (_N11935));
	// LUT = I0&~I1&~I2&I3&I4 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N537_4  */ #(
            .INIT(32'b00000000000100000000000000000000))
        \u_touch_top/u_touch_dri/N537_4  (
            .Z (_N11897),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [6] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [7] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [10] ),
            .I3 (\u_touch_top/u_touch_dri/cnt_time [15] ),
            .I4 (_N10457));
	// LUT = ~I0&~I1&I2&~I3&I4 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N537_5  */ #(
            .INIT(32'b00100000000000000000000000000000))
        \u_touch_top/u_touch_dri/N537_5  (
            .Z (\u_touch_top/u_touch_dri/N1629 [5] ),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [11] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [13] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [14] ),
            .I3 (_N11890),
            .I4 (_N11897));
	// LUT = I0&~I1&I2&I3&I4 ;

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N559[0]_1  */ #(
            .INIT(4'b0010))
        \u_touch_top/u_touch_dri/N559[0]_1  (
            .Z (\u_touch_top/u_touch_dri/N559 [0] ),
            .I0 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [0] ));
	// LUT = I0&~I1 ;
	// ../../rtl/touch/touch_dri.v:102

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N589_2  */ #(
            .INIT(16'b1011101000110000))
        \u_touch_top/u_touch_dri/N589_2  (
            .Z (_N11966),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I1 (\u_touch_top/u_touch_dri/st_done ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [0] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = (I0&I3)|(~I1&I2) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N592_or[0]_2  */ #(
            .INIT(32'b10101110000011001010101000000000))
        \u_touch_top/u_touch_dri/N592_or[0]_2  (
            .Z (_N11968),
            .I0 (\u_touch_top/u_touch_dri/N70 ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I2 (\u_touch_top/u_touch_dri/N1629 [5] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [0] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = (I1&~I2&I4)|(I0&I3) ;

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N614_2  */ #(
            .INIT(8'b10000000))
        \u_touch_top/u_touch_dri/N614_2  (
            .Z (\u_touch_top/u_touch_dri/N614 ),
            .I0 (\u_touch_top/once_byte_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [5] ));
	// LUT = I0&I1&I2 ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N641  */ #(
            .INIT(16'b1110000000000000))
        \u_touch_top/u_touch_dri/N641_vname  (
            .Z (\u_touch_top/u_touch_dri/N641 ),
            .I0 (\u_lcd_rgb_char/u_clk_div/N40 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [2] ));
    // defparam \u_touch_top/u_touch_dri/N641_vname .orig_name = \u_touch_top/u_touch_dri/N641 ;
	// LUT = (I1&I2&I3)|(I0&I2&I3) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N642  */ #(
            .INIT(32'b00000000000000001000100000100000))
        \u_touch_top/u_touch_dri/N642_vname  (
            .Z (\u_touch_top/u_touch_dri/N642 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I1 (\u_touch_top/u_touch_dri/st_done ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [2] ),
            .I3 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I4 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
    // defparam \u_touch_top/u_touch_dri/N642_vname .orig_name = \u_touch_top/u_touch_dri/N642 ;
	// LUT = (I0&~I1&I2&~I3&~I4)|(I0&I1&I3&~I4) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N647_1_9  */ #(
            .INIT(16'b0000000100000000))
        \u_touch_top/u_touch_dri/N647_1_9  (
            .Z (_N11956),
            .I0 (\u_touch_top/u_touch_dri/chip_version [2] ),
            .I1 (\u_touch_top/u_touch_dri/chip_version [3] ),
            .I2 (\u_touch_top/u_touch_dri/chip_version [4] ),
            .I3 (_N10246));
	// LUT = ~I0&~I1&~I2&I3 ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N647_1_11  */ #(
            .INIT(16'b0000000000000001))
        \u_touch_top/u_touch_dri/N647_1_11  (
            .Z (_N11958),
            .I0 (\u_touch_top/u_touch_dri/chip_version [9] ),
            .I1 (\u_touch_top/u_touch_dri/chip_version [10] ),
            .I2 (\u_touch_top/u_touch_dri/chip_version [11] ),
            .I3 (\u_touch_top/u_touch_dri/chip_version [14] ));
	// LUT = ~I0&~I1&~I2&~I3 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N647_1_13  */ #(
            .INIT(32'b00000000000000010000000000000000))
        \u_touch_top/u_touch_dri/N647_1_13  (
            .Z (_N11960),
            .I0 (\u_touch_top/u_touch_dri/chip_version [5] ),
            .I1 (\u_touch_top/u_touch_dri/chip_version [6] ),
            .I2 (\u_touch_top/u_touch_dri/chip_version [7] ),
            .I3 (\u_touch_top/u_touch_dri/chip_version [8] ),
            .I4 (_N11958));
	// LUT = ~I0&~I1&~I2&~I3&I4 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N666  */ #(
            .INIT(32'b00000000000000001000100000100000))
        \u_touch_top/u_touch_dri/N666_vname  (
            .Z (\u_touch_top/u_touch_dri/N666 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I1 (\u_touch_top/u_touch_dri/st_done ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [2] ),
            .I3 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I4 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
    // defparam \u_touch_top/u_touch_dri/N666_vname .orig_name = \u_touch_top/u_touch_dri/N666 ;
	// LUT = (I0&~I1&I2&~I3&~I4)|(I0&I1&I3&~I4) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N716  */ #(
            .INIT(16'b0100000000000000))
        \u_touch_top/u_touch_dri/N716_vname  (
            .Z (\u_touch_top/u_touch_dri/N716 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [5] ));
    // defparam \u_touch_top/u_touch_dri/N716_vname .orig_name = \u_touch_top/u_touch_dri/N716 ;
	// LUT = ~I0&I1&I2&I3 ;

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N739  */ #(
            .INIT(8'b10000000))
        \u_touch_top/u_touch_dri/N739_vname  (
            .Z (\u_touch_top/u_touch_dri/N739 ),
            .I0 (\u_touch_top/once_byte_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [5] ));
    // defparam \u_touch_top/u_touch_dri/N739_vname .orig_name = \u_touch_top/u_touch_dri/N739 ;
	// LUT = I0&I1&I2 ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N863_1  */ #(
            .INIT(4'b1110))
        \u_touch_top/u_touch_dri/N863_1  (
            .Z (\u_touch_top/u_touch_dri/N1281 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N863_6  */ #(
            .INIT(32'b11111111101010101111111110101000))
        \u_touch_top/u_touch_dri/N863_6  (
            .Z (\u_touch_top/u_touch_dri/N863 ),
            .I0 (\u_touch_top/once_byte_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I4 (\u_touch_top/u_touch_dri/N1281 ));
	// LUT = (I0&I4)|(I3)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N876_8  */ #(
            .INIT(32'b11111111111011001110110011101100))
        \u_touch_top/u_touch_dri/N876_8  (
            .Z (_N11923),
            .I0 (\u_touch_top/i2c_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I4 (\u_touch_top/u_touch_dri/N1629 [5] ));
	// LUT = (I3&I4)|(I0&I2)|(I1) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N891_0_3  */ #(
            .INIT(16'b1111111111111110))
        \u_touch_top/u_touch_dri/N891_0_3  (
            .Z (\u_touch_top/u_touch_dri/N1201 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ));
	// LUT = (I3)|(I2)|(I1)|(I0) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N891_1_2  */ #(
            .INIT(16'b1010101010101000))
        \u_touch_top/u_touch_dri/N891_1_2  (
            .Z (_N11925),
            .I0 (\u_touch_top/i2c_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [7] ));
	// LUT = (I0&I3)|(I0&I2)|(I0&I1) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N905_2  */ #(
            .INIT(32'b11111111111111111110110010100000))
        \u_touch_top/u_touch_dri/N905_2  (
            .Z (_N11928),
            .I0 (\u_touch_top/i2c_done ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I4 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ));
	// LUT = (I4)|(I1&I3)|(I0&I2) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N905_5  */ #(
            .INIT(32'b11111111111111111111111011111010))
        \u_touch_top/u_touch_dri/N905_5  (
            .Z (\u_touch_top/u_touch_dri/N905 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I2 (\u_touch_top/u_touch_dri/N1281 ),
            .I3 (_N10532),
            .I4 (_N11928));
	// LUT = (I4)|(I1&I3)|(I2)|(I0) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N924  */ #(
            .INIT(32'b00000000000000001000100000100000))
        \u_touch_top/u_touch_dri/N924_vname  (
            .Z (\u_touch_top/u_touch_dri/N924 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I1 (\u_touch_top/u_touch_dri/st_done ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [2] ),
            .I3 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I4 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
    // defparam \u_touch_top/u_touch_dri/N924_vname .orig_name = \u_touch_top/u_touch_dri/N924 ;
	// LUT = (I0&~I1&I2&~I3&~I4)|(I0&I1&I3&~I4) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N933  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_touch_dri/N933_vname  (
            .Z (\u_touch_top/u_touch_dri/N933 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I1 (\u_touch_top/u_touch_dri/next_state [3] ));
    // defparam \u_touch_top/u_touch_dri/N933_vname .orig_name = \u_touch_top/u_touch_dri/N933 ;
	// LUT = I0&I1 ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N935  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_touch_dri/N935_vname  (
            .Z (\u_touch_top/u_touch_dri/N935 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ),
            .I1 (\u_touch_top/u_touch_dri/next_state [3] ));
    // defparam \u_touch_top/u_touch_dri/N935_vname .orig_name = \u_touch_top/u_touch_dri/N935 ;
	// LUT = I0&I1 ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N937  */ #(
            .INIT(32'b00000000000000000000011100000000))
        \u_touch_top/u_touch_dri/N937_vname  (
            .Z (\u_touch_top/u_touch_dri/N937 ),
            .I0 (\u_touch_top/i2c_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .I2 (\u_touch_top/u_touch_dri/N1201 ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (_N11925));
    // defparam \u_touch_top/u_touch_dri/N937_vname .orig_name = \u_touch_top/u_touch_dri/N937 ;
	// LUT = (~I1&~I2&I3&~I4)|(~I0&~I2&I3&~I4) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N944  */ #(
            .INIT(32'b00000000000000000000011100000000))
        \u_touch_top/u_touch_dri/N944_vname  (
            .Z (\u_touch_top/u_touch_dri/N944 ),
            .I0 (\u_touch_top/i2c_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I2 (\u_touch_top/u_touch_dri/N1281 ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I4 (_N11923));
    // defparam \u_touch_top/u_touch_dri/N944_vname .orig_name = \u_touch_top/u_touch_dri/N944 ;
	// LUT = (~I1&~I2&I3&~I4)|(~I0&~I2&I3&~I4) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N945  */ #(
            .INIT(4'b1000))
        \u_touch_top/u_touch_dri/N945_vname  (
            .Z (\u_touch_top/u_touch_dri/N945 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I1 (\u_touch_top/u_touch_dri/next_state [5] ));
    // defparam \u_touch_top/u_touch_dri/N945_vname .orig_name = \u_touch_top/u_touch_dri/N945 ;
	// LUT = I0&I1 ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N948  */ #(
            .INIT(8'b10000000))
        \u_touch_top/u_touch_dri/N948_vname  (
            .Z (\u_touch_top/u_touch_dri/N948 ),
            .I0 (\u_touch_top/once_byte_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [5] ));
    // defparam \u_touch_top/u_touch_dri/N948_vname .orig_name = \u_touch_top/u_touch_dri/N948 ;
	// LUT = I0&I1&I2 ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT5M /* \u_touch_top/u_touch_dri/N951_2  */ #(
            .INIT(32'b01010101010101010000000000000001))
        \u_touch_top/u_touch_dri/N951_2  (
            .Z (_N11940),
            .I0 (\u_touch_top/u_touch_dri/N474 ),
            .I1 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [5] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [1] ),
            .ID (\u_touch_top/u_touch_dri/next_state [2] ));
	// LUT = (~ID&~I1&~I2&~I3&~I4)|(~I0&I4) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N951_7  */ #(
            .INIT(32'b11111111111111111111110111111100))
        \u_touch_top/u_touch_dri/N951_7  (
            .Z (_N11945),
            .I0 (\u_touch_top/u_touch_dri/N863 ),
            .I1 (\u_touch_top/u_touch_dri/N944 ),
            .I2 (\u_touch_top/u_touch_dri/next_state [0] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [5] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [6] ));
	// LUT = (I4)|(~I0&I3)|(I2)|(I1) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N961  */ #(
            .INIT(32'b00000000000000000000000000100011))
        \u_touch_top/u_touch_dri/N961_vname  (
            .Z (\u_touch_top/u_touch_dri/N961 ),
            .I0 (\u_touch_top/u_touch_dri/N905 ),
            .I1 (\u_touch_top/u_touch_dri/N937 ),
            .I2 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I3 (_N11940),
            .I4 (_N11945));
    // defparam \u_touch_top/u_touch_dri/N961_vname .orig_name = \u_touch_top/u_touch_dri/N961 ;
	// LUT = (~I1&~I2&~I3&~I4)|(I0&~I1&~I3&~I4) ;

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N1074  */ #(
            .INIT(8'b11100000))
        \u_touch_top/u_touch_dri/N1074_vname  (
            .Z (\u_touch_top/u_touch_dri/N1074 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [2] ));
    // defparam \u_touch_top/u_touch_dri/N1074_vname .orig_name = \u_touch_top/u_touch_dri/N1074 ;
	// LUT = (I1&I2)|(I0&I2) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1206  */ #(
            .INIT(32'b11111111111111100000000000000000))
        \u_touch_top/u_touch_dri/N1206_vname  (
            .Z (\u_touch_top/u_touch_dri/N1206 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [3] ));
    // defparam \u_touch_top/u_touch_dri/N1206_vname .orig_name = \u_touch_top/u_touch_dri/N1206 ;
	// LUT = (I3&I4)|(I2&I4)|(I1&I4)|(I0&I4) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT5M /* \u_touch_top/u_touch_dri/N1218  */ #(
            .INIT(32'b00000101000001010000111100011111))
        \u_touch_top/u_touch_dri/N1218_vname  (
            .Z (\u_touch_top/u_touch_dri/N1218 ),
            .I0 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I4 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .ID (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ));
    // defparam \u_touch_top/u_touch_dri/N1218_vname .orig_name = \u_touch_top/u_touch_dri/N1218 ;
	// LUT = (~ID&~I1&~I3&~I4)|(~I2&~I4)|(~I0&~I2) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1297_4  */ #(
            .INIT(32'b11111111111111111111111011110000))
        \u_touch_top/u_touch_dri/N1297_4  (
            .Z (\u_touch_top/u_touch_dri/N1297 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I2 (\u_touch_top/u_touch_dri/N1300 [5] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (_N10481));
	// LUT = (I4)|(I1&I3)|(I0&I3)|(I2) ;

    GTP_LUT3 /* \u_touch_top/u_touch_dri/N1300_and[4][6]  */ #(
            .INIT(8'b10000000))
        \u_touch_top/u_touch_dri/N1300_and[4][6]  (
            .Z (\u_touch_top/u_touch_dri/N1300 [4] ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I1 (\u_touch_top/u_touch_dri/coord_reg [4] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [5] ));
	// LUT = I0&I1&I2 ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N1300_and[6]_1  */ #(
            .INIT(16'b1110101011000000))
        \u_touch_top/u_touch_dri/N1300_and[6]_1  (
            .Z (\u_touch_top/u_touch_dri/N1300 [5] ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ));
	// LUT = (I0&I3)|(I1&I2) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1300_inv[6]  */ #(
            .INIT(32'b00010001010101010001001101011111))
        \u_touch_top/u_touch_dri/N1300_inv[6]  (
            .Z (\u_touch_top/u_touch_dri/N1300 [7] ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I1 (\u_touch_top/u_touch_dri/N1281 ),
            .I2 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [5] ));
	// LUT = (~I2&~I3&~I4)|(~I1&~I2&~I4)|(~I0&~I3)|(~I0&~I1) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1300_or[0]  */ #(
            .INIT(32'b11101010110000001010101000000000))
        \u_touch_top/u_touch_dri/N1300_or[0]  (
            .Z (\u_touch_top/u_touch_dri/N1300 [0] ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I2 (\u_touch_top/u_touch_dri/coord_reg [0] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [5] ));
	// LUT = (I1&I2&I4)|(I0&I3) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1300_or[1]  */ #(
            .INIT(32'b11101100101000001010000010100000))
        \u_touch_top/u_touch_dri/N1300_or[1]  (
            .Z (\u_touch_top/u_touch_dri/N1300 [1] ),
            .I0 (\u_touch_top/u_touch_dri/N945 ),
            .I1 (\u_touch_top/u_touch_dri/N1281 ),
            .I2 (\u_touch_top/u_touch_dri/coord_reg [0] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I4 (\u_touch_top/u_touch_dri/touch_s_reg [1] ));
	// LUT = (I1&I3&I4)|(I0&I2) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1300_or[2]  */ #(
            .INIT(32'b11101010110000001010101000000000))
        \u_touch_top/u_touch_dri/N1300_or[2]  (
            .Z (\u_touch_top/u_touch_dri/N1300 [2] ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I1 (\u_touch_top/u_touch_dri/N1281 ),
            .I2 (\u_touch_top/u_touch_dri/coord_reg [4] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = (I1&I2&I4)|(I0&I3) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1300_or[3]  */ #(
            .INIT(32'b11101010110000001010101000000000))
        \u_touch_top/u_touch_dri/N1300_or[3]  (
            .Z (\u_touch_top/u_touch_dri/N1300 [3] ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ),
            .I1 (\u_touch_top/u_touch_dri/N1281 ),
            .I2 (\u_touch_top/u_touch_dri/coord_reg [4] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = (I1&I2&I4)|(I0&I3) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1300_or[5]  */ #(
            .INIT(32'b11111110000000001111000000000000))
        \u_touch_top/u_touch_dri/N1300_or[5]  (
            .Z (\u_touch_top/u_touch_dri/N1300 [6] ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I2 (\u_touch_top/u_touch_dri/N945 ),
            .I3 (\u_touch_top/u_touch_dri/coord_reg [4] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = (I1&I3&I4)|(I0&I3&I4)|(I2&I3) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1345_1  */ #(
            .INIT(32'b11101110101010101110110010100000))
        \u_touch_top/u_touch_dri/N1345_1  (
            .Z (_N10481),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I1 (\u_touch_top/u_touch_dri/N1281 ),
            .I2 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [5] ));
	// LUT = (I0&I4)|(I1&I3)|(I0&I2) ;

    GTP_LUT5M /* \u_touch_top/u_touch_dri/N1450_1  */ #(
            .INIT(32'b11111010111110101111000011100000))
        \u_touch_top/u_touch_dri/N1450_1  (
            .Z (\u_touch_top/u_touch_dri/N1216 ),
            .I0 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I4 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .ID (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ));
	// LUT = (I2&I4)|(I0&I4)|(I2&I3)|(I1&I2)|(ID&I2) ;

    GTP_LUT5M /* \u_touch_top/u_touch_dri/N1450_5  */ #(
            .INIT(32'b11111111111111101111111011111100))
        \u_touch_top/u_touch_dri/N1450_5  (
            .Z (\u_touch_top/u_touch_dri/N1450 ),
            .I0 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I1 (\u_touch_top/u_touch_dri/N1206 ),
            .I2 (\u_touch_top/u_touch_dri/N945 ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I4 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .ID (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ));
	// LUT = (I3&I4)|(I0&I4)|(ID&I3)|(I2)|(I1) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N1453  */ #(
            .INIT(16'b1111111011110000))
        \u_touch_top/u_touch_dri/N1453_vname  (
            .Z (\u_touch_top/u_touch_dri/N1453 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I2 (\u_touch_top/u_touch_dri/N1206 ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ));
    // defparam \u_touch_top/u_touch_dri/N1453_vname .orig_name = \u_touch_top/u_touch_dri/N1453 ;
	// LUT = (I1&I3)|(I0&I3)|(I2) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N1491_4  */ #(
            .INIT(16'b0001000000000000))
        \u_touch_top/u_touch_dri/N1491_4  (
            .Z (_N10560),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [11] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [12] ),
            .I2 (_N10518),
            .I3 (_N10519));
	// LUT = ~I0&~I1&I2&I3 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1492_6  */ #(
            .INIT(32'b10000000000000000000000000000000))
        \u_touch_top/u_touch_dri/N1492_6  (
            .Z (_N12199),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [4] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [8] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [10] ),
            .I3 (_N10517),
            .I4 (_N10560));
	// LUT = I0&I1&I2&I3&I4 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1494  */ #(
            .INIT(32'b11001100100010001100010000000000))
        \u_touch_top/u_touch_dri/N1494_vname  (
            .Z (\u_touch_top/u_touch_dri/N1494 ),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [13] ),
            .I1 (\u_touch_top/u_touch_dri/next_state [1] ),
            .I2 (_N574),
            .I3 (_N10519),
            .I4 (_N12199));
    // defparam \u_touch_top/u_touch_dri/N1494_vname .orig_name = \u_touch_top/u_touch_dri/N1494 ;
	// LUT = (I0&I1&I4)|(I1&I2&I3)|(~I0&I1&I3) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT4 /* \u_touch_top/u_touch_dri/N1497  */ #(
            .INIT(16'b0011101111111111))
        \u_touch_top/u_touch_dri/N1497_vname  (
            .Z (\u_touch_top/u_touch_dri/N1497 ),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [13] ),
            .I1 (\u_touch_top/u_touch_dri/next_state [1] ),
            .I2 (_N574),
            .I3 (_N10519));
    // defparam \u_touch_top/u_touch_dri/N1497_vname .orig_name = \u_touch_top/u_touch_dri/N1497 ;
	// LUT = (~I3)|(I0&~I2)|(~I1) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1529  */ #(
            .INIT(32'b11111000000000000000000000000000))
        \u_touch_top/u_touch_dri/N1529_vname  (
            .Z (\u_touch_top/u_touch_dri/N1529 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [2] ));
    // defparam \u_touch_top/u_touch_dri/N1529_vname .orig_name = \u_touch_top/u_touch_dri/N1529 ;
	// LUT = (I2&I3&I4)|(I0&I1&I3&I4) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1569  */ #(
            .INIT(32'b11111000000000001000100000000000))
        \u_touch_top/u_touch_dri/N1569_vname  (
            .Z (\u_touch_top/u_touch_dri/N1569 ),
            .I0 (\u_touch_top/i2c_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I4 (_N10532));
    // defparam \u_touch_top/u_touch_dri/N1569_vname .orig_name = \u_touch_top/u_touch_dri/N1569 ;
	// LUT = (I2&I3&I4)|(I0&I1&I3) ;
	// ../../rtl/touch/touch_dri.v:214

    GTP_LUT2 /* \u_touch_top/u_touch_dri/N1610_2  */ #(
            .INIT(4'b1110))
        \u_touch_top/u_touch_dri/N1610_2  (
            .Z (_N11905),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ));
	// LUT = (I1)|(I0) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/N1610_3  */ #(
            .INIT(32'b11111111111111111111111111111110))
        \u_touch_top/u_touch_dri/N1610_3  (
            .Z (\u_touch_top/u_touch_dri/N1610 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [7] ),
            .I4 (_N11905));
	// LUT = (I4)|(I3)|(I2)|(I1)|(I0) ;

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/bit_ctrl  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/bit_ctrl  (
            .Q (\u_touch_top/bit_ctrl ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1074 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9402));
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT2 /* \u_touch_top/u_touch_dri/bit_ctrl_0  */ #(
            .INIT(4'b1110))
        \u_touch_top/u_touch_dri/bit_ctrl_0  (
            .Z (_N9403),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I1 (\u_touch_top/u_touch_dri/ft_flag ));
	// LUT = (I1)|(I0) ;

    GTP_LUT2 /* \u_touch_top/u_touch_dri/bit_ctrl_32  */ #(
            .INIT(4'b0001))
        \u_touch_top/u_touch_dri/bit_ctrl_32  (
            .Z (_N9402),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I1 (\u_touch_top/u_touch_dri/ft_flag ));
	// LUT = ~I0&~I1 ;

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[0]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1569 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9426));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[1]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1569 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9468));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[2]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1569 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9512));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[3]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1569 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9551));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[4]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1569 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9596));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[5]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1569 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9641));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[6]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1569 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9679));
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[7:0]_0  */ #(
            .INIT(16'b1101000011110000))
        \u_touch_top/u_touch_dri/chip_version[7:0]_0  (
            .Z (_N9426),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/i2c_data_r [0] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ));
	// LUT = (I2&~I3)|(I1&I2)|(~I0&I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[7:0]_3  */ #(
            .INIT(16'b1101000011110000))
        \u_touch_top/u_touch_dri/chip_version[7:0]_3  (
            .Z (_N9468),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/i2c_data_r [1] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ));
	// LUT = (I2&~I3)|(I1&I2)|(~I0&I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[7:0]_6  */ #(
            .INIT(16'b1111001011110000))
        \u_touch_top/u_touch_dri/chip_version[7:0]_6  (
            .Z (_N9512),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/i2c_data_r [2] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ));
	// LUT = (I0&~I1&I3)|(I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[7:0]_9  */ #(
            .INIT(16'b1101000011110000))
        \u_touch_top/u_touch_dri/chip_version[7:0]_9  (
            .Z (_N9551),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/i2c_data_r [3] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ));
	// LUT = (I2&~I3)|(I1&I2)|(~I0&I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[7:0]_79  */ #(
            .INIT(16'b1111001011110000))
        \u_touch_top/u_touch_dri/chip_version[7:0]_79  (
            .Z (_N9596),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/i2c_data_r [4] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ));
	// LUT = (I0&~I1&I3)|(I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[7:0]_117  */ #(
            .INIT(16'b1101000011110000))
        \u_touch_top/u_touch_dri/chip_version[7:0]_117  (
            .Z (_N9641),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/i2c_data_r [5] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ));
	// LUT = (I2&~I3)|(I1&I2)|(~I0&I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[7:0]_151  */ #(
            .INIT(16'b1111001011110000))
        \u_touch_top/u_touch_dri/chip_version[7:0]_151  (
            .Z (_N9679),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/i2c_data_r [6] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ));
	// LUT = (I0&~I1&I3)|(I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[7:0]_189  */ #(
            .INIT(16'b1101000011110000))
        \u_touch_top/u_touch_dri/chip_version[7:0]_189  (
            .Z (_N9724),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/i2c_data_r [7] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ));
	// LUT = (I2&~I3)|(I1&I2)|(~I0&I2) ;

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[7]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1569 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9724));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[8]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1529 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9759));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[9]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1529 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9791));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[10]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1529 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9827));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[11]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1529 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9859));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[12]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [12] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1529 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9907));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[13]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [13] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1529 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9955));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[14]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [14] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1529 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N10009));
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[15:8]_0  */ #(
            .INIT(16'b1111111100001000))
        \u_touch_top/u_touch_dri/chip_version[15:8]_0  (
            .Z (_N9759),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/i2c_data_r [0] ));
	// LUT = (I3)|(I0&I1&~I2) ;

    GTP_LUT3 /* \u_touch_top/u_touch_dri/chip_version[15:8]_2  */ #(
            .INIT(8'b00010000))
        \u_touch_top/u_touch_dri/chip_version[15:8]_2  (
            .Z (_N10519),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [14] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [15] ),
            .I2 (_N10457));
	// LUT = ~I0&~I1&I2 ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[15:8]_3  */ #(
            .INIT(16'b1111111100001000))
        \u_touch_top/u_touch_dri/chip_version[15:8]_3  (
            .Z (_N9791),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/i2c_data_r [1] ));
	// LUT = (I3)|(I0&I1&~I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[15:8]_6  */ #(
            .INIT(16'b1111111100001000))
        \u_touch_top/u_touch_dri/chip_version[15:8]_6  (
            .Z (_N9827),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/i2c_data_r [2] ));
	// LUT = (I3)|(I0&I1&~I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[15:8]_88  */ #(
            .INIT(16'b1111011100000000))
        \u_touch_top/u_touch_dri/chip_version[15:8]_88  (
            .Z (_N9859),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/i2c_data_r [3] ));
	// LUT = (I2&I3)|(~I1&I3)|(~I0&I3) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[15:8]_101  */ #(
            .INIT(16'b1111011100000000))
        \u_touch_top/u_touch_dri/chip_version[15:8]_101  (
            .Z (_N9907),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/i2c_data_r [4] ));
	// LUT = (I2&I3)|(~I1&I3)|(~I0&I3) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[15:8]_114  */ #(
            .INIT(16'b1111011100000000))
        \u_touch_top/u_touch_dri/chip_version[15:8]_114  (
            .Z (_N9955),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/i2c_data_r [5] ));
	// LUT = (I2&I3)|(~I1&I3)|(~I0&I3) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[15:8]_131  */ #(
            .INIT(16'b1111011100000000))
        \u_touch_top/u_touch_dri/chip_version[15:8]_131  (
            .Z (_N10046),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/i2c_data_r [7] ));
	// LUT = (I2&I3)|(~I1&I3)|(~I0&I3) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/chip_version[15:8]_149  */ #(
            .INIT(16'b1111111100001000))
        \u_touch_top/u_touch_dri/chip_version[15:8]_149  (
            .Z (_N10009),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/i2c_data_r [6] ));
	// LUT = (I3)|(I0&I1&~I2) ;

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/chip_version[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/chip_version[15]  (
            .Q (\u_touch_top/u_touch_dri/chip_version [15] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1529 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N10046));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[0]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [0] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[1]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [1] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[2]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [2] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[3]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [3] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[4]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [4] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[5]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [5] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[6]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [6] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[7]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [7] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[8]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [8] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[9]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [9] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[10]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [10] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[11]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [11] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[12]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [12] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [12] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[13]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [13] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [13] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[14]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [14] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [14] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[15]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [15] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [15] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[16]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[16]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [16] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [16] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[17]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[17]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [17] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [17] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[18]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[18]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [18] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [18] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_C /* \u_touch_top/u_touch_dri/cnt_time[19]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time[19]  (
            .Q (\u_touch_top/u_touch_dri/cnt_time [19] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N559 [19] ));
	// ../../rtl/touch/touch_dri.v:102

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/cnt_time_en  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cnt_time_en_vname  (
            .Q (\u_touch_top/u_touch_dri/cnt_time_en ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (1'b1),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N11807));
    // defparam \u_touch_top/u_touch_dri/cnt_time_en_vname .orig_name = \u_touch_top/u_touch_dri/cnt_time_en ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5 /* \u_touch_top/u_touch_dri/cnt_time_en_ce_mux  */ #(
            .INIT(32'b11111111111111000101000001011100))
        \u_touch_top/u_touch_dri/cnt_time_en_ce_mux  (
            .Z (_N11807),
            .I0 (\u_touch_top/u_touch_dri/N474 ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time_en ),
            .I2 (\u_touch_top/u_touch_dri/next_state [1] ),
            .I3 (_N11966),
            .I4 (_N11968));
	// LUT = (I3&I4)|(I2&I4)|(I1&~I2&~I3)|(~I0&I2) ;

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/coord_reg[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/coord_reg[0]  (
            .Q (\u_touch_top/u_touch_dri/coord_reg [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N666 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/ft_flag ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/coord_reg[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/coord_reg[4]  (
            .Q (\u_touch_top/u_touch_dri/coord_reg [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N666 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N166 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT2 /* \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_1  */ #(
            .INIT(4'b0100))
        \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_1  (
            .Z (\u_touch_top/u_touch_dri/next_state [0] ),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
	// LUT = ~I0&I1 ;
	// ../../rtl/touch/touch_dri.v:124

    GTP_LUT3 /* \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_4  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_4  (
            .Z (\u_touch_top/u_touch_dri/_N48 ),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:124

    GTP_LUT3 /* \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_7  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_7  (
            .Z (\u_touch_top/u_touch_dri/_N51 ),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [2] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [1] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:124

    GTP_LUT4 /* \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_11  */ #(
            .INIT(16'b1011100000110000))
        \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_11  (
            .Z (\u_touch_top/u_touch_dri/_N55 ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/st_done ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [3] ),
            .I3 (\u_touch_top/u_touch_dri/cur_state_reg [2] ));
	// LUT = (I0&I1&I3)|(~I1&I2) ;
	// ../../rtl/touch/touch_dri.v:124

    GTP_LUT3 /* \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_20  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_20  (
            .Z (\u_touch_top/u_touch_dri/_N64 ),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [5] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [4] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:124

    GTP_LUT3 /* \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_23  */ #(
            .INIT(8'b11100100))
        \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_23  (
            .Z (\u_touch_top/u_touch_dri/_N67 ),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [6] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [5] ));
	// LUT = (I0&I2)|(~I0&I1) ;
	// ../../rtl/touch/touch_dri.v:124

    GTP_LUT5M /* \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_24_3  */ #(
            .INIT(32'b11111101111111001010101010101010))
        \u_touch_top/u_touch_dri/cur_state_fsm[6:0]_24_3  (
            .Z (\u_touch_top/u_touch_dri/_N61 ),
            .I0 (\u_touch_top/u_touch_dri/ft_flag ),
            .I1 (\u_touch_top/u_touch_dri/cur_state_reg [6] ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [3] ),
            .I3 (\u_touch_top/u_touch_dri/cur_state_reg [2] ),
            .I4 (\u_touch_top/u_touch_dri/st_done ),
            .ID (\u_touch_top/u_touch_dri/cur_state_reg [4] ));
	// LUT = (ID&~I4)|(~I0&I3&I4)|(I2&I4)|(I1&I4) ;

(* syn_encoding="onehot" *)    GTP_DFF_P /* \u_touch_top/u_touch_dri/cur_state_reg[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b1))
        \u_touch_top/u_touch_dri/cur_state_reg[0]  (
            .Q (\u_touch_top/u_touch_dri/cur_state_reg [0] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/next_state [0] ),
            .P (\u_lcd_rgb_char/u_binary2bcd_x/N0 ));
	// ../../rtl/touch/touch_dri.v:124

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_touch_dri/cur_state_reg[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cur_state_reg[1]  (
            .Q (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N48 ));
	// ../../rtl/touch/touch_dri.v:124

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_touch_dri/cur_state_reg[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cur_state_reg[2]  (
            .Q (\u_touch_top/u_touch_dri/cur_state_reg [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N51 ));
	// ../../rtl/touch/touch_dri.v:124

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_touch_dri/cur_state_reg[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cur_state_reg[3]  (
            .Q (\u_touch_top/u_touch_dri/cur_state_reg [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N55 ));
	// ../../rtl/touch/touch_dri.v:124

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_touch_dri/cur_state_reg[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cur_state_reg[4]  (
            .Q (\u_touch_top/u_touch_dri/cur_state_reg [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N61 ));
	// ../../rtl/touch/touch_dri.v:124

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_touch_dri/cur_state_reg[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cur_state_reg[5]  (
            .Q (\u_touch_top/u_touch_dri/cur_state_reg [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N64 ));
	// ../../rtl/touch/touch_dri.v:124

(* syn_encoding="onehot" *)    GTP_DFF_C /* \u_touch_top/u_touch_dri/cur_state_reg[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/cur_state_reg[6]  (
            .Q (\u_touch_top/u_touch_dri/cur_state_reg [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N67 ));
	// ../../rtl/touch/touch_dri.v:124

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[0]  (
            .Q (data[0]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [0] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[1]  (
            .Q (data[1]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [1] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[2]  (
            .Q (data[2]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [2] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[3]  (
            .Q (data[3]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [3] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[4]  (
            .Q (data[4]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [4] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[5]  (
            .Q (data[5]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [5] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[6]  (
            .Q (data[6]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [6] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[7]  (
            .Q (data[7]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [7] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[8]  (
            .Q (data[8]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [8] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[9]  (
            .Q (data[9]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [9] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[10]  (
            .Q (data[10]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [10] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[11]  (
            .Q (data[11]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [11] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[12]  (
            .Q (data[12]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [12] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[13]  (
            .Q (data[13]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [13] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[14]  (
            .Q (data[14]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [14] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[15]  (
            .Q (data[15]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_y_coord [15] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[16]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[16]  (
            .Q (data[16]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [0] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[17]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[17]  (
            .Q (data[17]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [1] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[18]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[18]  (
            .Q (data[18]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [2] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[19]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[19]  (
            .Q (data[19]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [3] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[20]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[20]  (
            .Q (data[20]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [4] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[21]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[21]  (
            .Q (data[21]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [5] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[22]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[22]  (
            .Q (data[22]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [6] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[23]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[23]  (
            .Q (data[23]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [7] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[24]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[24]  (
            .Q (data[24]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [8] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[25]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[25]  (
            .Q (data[25]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [9] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[26]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[26]  (
            .Q (data[26]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [10] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[27]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[27]  (
            .Q (data[27]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [11] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[28]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[28]  (
            .Q (data[28]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [12] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[29]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[29]  (
            .Q (data[29]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [13] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[30]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[30]  (
            .Q (data[30]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [14] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/data[31]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/data[31]  (
            .Q (data[31]),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/touch_valid ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/tp_x_coord [15] ));
	// ../../rtl/touch/touch_dri.v:113

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_3  */ #(
            .INIT(32'b10101000101000001000100000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_3  (
            .Z (\u_touch_top/u_touch_dri/_N70 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [5] ));
	// LUT = (I0&I2&I4)|(I0&I1&I3) ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT3 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_7  */ #(
            .INIT(8'b01000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_7  (
            .Z (\u_touch_top/u_touch_dri/_N74 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = ~I0&I1&I2 ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT4 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_14  */ #(
            .INIT(16'b0100000000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_14  (
            .Z (\u_touch_top/u_touch_dri/_N81 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I3 (\u_touch_top/u_touch_dri/flow_cnt_reg [7] ));
	// LUT = ~I0&I1&I2&I3 ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_18_3  */ #(
            .INIT(32'b11101110101010101110110010100000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_18_3  (
            .Z (_N11990),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I3 (\u_touch_top/u_touch_dri/_N70 ),
            .I4 (\u_touch_top/u_touch_dri/_N74 ));
	// LUT = (I0&I4)|(I1&I3)|(I0&I2) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_18_5  */ #(
            .INIT(32'b11111111111111111111111111101100))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_18_5  (
            .Z (\u_touch_top/u_touch_dri/_N85 ),
            .I0 (\u_touch_top/u_touch_dri/N474 ),
            .I1 (\u_touch_top/u_touch_dri/N614 ),
            .I2 (\u_touch_top/u_touch_dri/next_state [1] ),
            .I3 (\u_touch_top/u_touch_dri/_N81 ),
            .I4 (_N11990));
	// LUT = (I4)|(I3)|(I0&I2)|(I1) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_21_2  */ #(
            .INIT(32'b11111111111111111111111100010000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_21_2  (
            .Z (_N11899),
            .I0 (\u_lcd_rgb_char/u_clk_div/N40 ),
            .I1 (\u_lcd_rgb_char/u_lcd_driver/h_sync [3] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [5] ));
	// LUT = (I4)|(I3)|(~I0&~I1&I2) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_24  */ #(
            .INIT(16'b1000000000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_24  (
            .Z (\u_touch_top/u_touch_dri/_N91 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = I0&I1&I2&I3 ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_28_2  */ #(
            .INIT(32'b11111111101010101111111110000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_28_2  (
            .Z (\u_touch_top/u_touch_dri/_N95 ),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I1 (\u_touch_top/u_touch_dri/N1629 [5] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I3 (\u_touch_top/u_touch_dri/_N91 ),
            .I4 (_N11899));
	// LUT = (I0&I4)|(I3)|(I0&I1&I2) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_31_2  */ #(
            .INIT(32'b11111111111111111111010011110000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_31_2  (
            .Z (_N11882),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = (I4)|(~I0&I1&I3)|(I2) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_32  */ #(
            .INIT(32'b11110000111100000100000000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_32  (
            .Z (\u_touch_top/u_touch_dri/_N99 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/once_byte_done ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [5] ),
            .I4 (_N11882));
	// LUT = (I2&I4)|(~I0&I1&I2&I3) ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_35  */ #(
            .INIT(32'b11111111111111111000000000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_35  (
            .Z (\u_touch_top/u_touch_dri/_N102 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (\u_touch_top/u_touch_dri/_N99 ));
	// LUT = (I4)|(I0&I1&I2&I3) ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_39_2  */ #(
            .INIT(32'b11110100111100000100010000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_39_2  (
            .Z (_N11901),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [5] ));
	// LUT = (I2&I4)|(~I0&I1&I3) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_40  */ #(
            .INIT(32'b11001100110011001100110010000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_40  (
            .Z (\u_touch_top/u_touch_dri/_N107 ),
            .I0 (\u_touch_top/once_byte_done ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (_N11901));
	// LUT = (I1&I4)|(I1&I3)|(I0&I1&I2) ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_44_2  */ #(
            .INIT(32'b11110100111100000100010000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_44_2  (
            .Z (_N11914),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/once_byte_done ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [5] ));
	// LUT = (I2&I4)|(~I0&I1&I3) ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_44_4  */ #(
            .INIT(16'b1111111111111000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_44_4  (
            .Z (\u_touch_top/u_touch_dri/_N111 ),
            .I0 (\u_touch_top/i2c_done ),
            .I1 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I3 (_N11914));
	// LUT = (I3)|(I2)|(I0&I1) ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_52  */ #(
            .INIT(32'b10000000100000001000000000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_52  (
            .Z (\u_touch_top/u_touch_dri/_N119 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = (I0&I1&I2&I4)|(I0&I1&I2&I3) ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5M /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_53_3  */ #(
            .INIT(32'b11111110111110101111100011110000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_53_3  (
            .Z (\u_touch_top/u_touch_dri/_N120 ),
            .I0 (\u_touch_top/u_touch_dri/_N111 ),
            .I1 (\u_touch_top/u_touch_dri/next_state [2] ),
            .I2 (\u_touch_top/u_touch_dri/_N119 ),
            .I3 (_N10532),
            .I4 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .ID (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ));
	// LUT = (I1&I3&I4)|(I0&I4)|(ID&I1&I3)|(I2) ;

    GTP_LUT5M /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_59  */ #(
            .INIT(32'b11101100111011001100110010001000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_59  (
            .Z (\u_touch_top/u_touch_dri/_N126 ),
            .I0 (\u_touch_top/u_touch_dri/N1629 [9] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I4 (\u_touch_top/u_touch_dri/next_state [2] ),
            .ID (\u_touch_top/u_touch_dri/next_state [3] ));
	// LUT = (I0&I2&I4)|(I1&I4)|(I1&I3)|(ID&I1) ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_64  */ #(
            .INIT(32'b11001000000000000100000000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_64  (
            .Z (\u_touch_top/u_touch_dri/_N131 ),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/i2c_done ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I4 (\u_touch_top/u_touch_dri/flow_cnt_reg [7] ));
	// LUT = (I0&I1&I3&I4)|(~I0&I1&I2&I3) ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT3 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_95  */ #(
            .INIT(8'b00000001))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_95  (
            .Z (_N10518),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [5] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [6] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [7] ));
	// LUT = ~I0&~I1&~I2 ;

    GTP_LUT2 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_96  */ #(
            .INIT(4'b0001))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_96  (
            .Z (_N10520),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [4] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [8] ));
	// LUT = ~I0&~I1 ;

    GTP_LUT4 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_97  */ #(
            .INIT(16'b0000000000000001))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_97  (
            .Z (_N10521),
            .I0 (\u_touch_top/u_touch_dri/next_state [3] ),
            .I1 (\u_touch_top/u_touch_dri/next_state [4] ),
            .I2 (\u_touch_top/u_touch_dri/next_state [5] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [6] ));
	// LUT = ~I0&~I1&~I2&~I3 ;

    GTP_LUT3 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_99  */ #(
            .INIT(8'b01000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_99  (
            .Z (_N10558),
            .I0 (\u_touch_top/i2c_ack ),
            .I1 (\u_touch_top/u_i2c_dri/cur_state_reg [3] ),
            .I2 (\u_touch_top/u_i2c_dri/st_done ));
	// LUT = ~I0&I1&I2 ;

    GTP_LUT5 /* \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_106  */ #(
            .INIT(32'b00000000000000010000000000000000))
        \u_touch_top/u_touch_dri/flow_cnt_fsm[3:0]_106  (
            .Z (_N10517),
            .I0 (\u_touch_top/u_touch_dri/cnt_time [0] ),
            .I1 (\u_touch_top/u_touch_dri/cnt_time [1] ),
            .I2 (\u_touch_top/u_touch_dri/cnt_time [2] ),
            .I3 (\u_touch_top/u_touch_dri/cnt_time [3] ),
            .I4 (\u_touch_top/u_touch_dri/cnt_time [9] ));
	// LUT = ~I0&~I1&~I2&~I3&I4 ;

(* syn_encoding="onehot" *)    GTP_DFF_PE /* \u_touch_top/u_touch_dri/flow_cnt_reg[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b1))
        \u_touch_top/u_touch_dri/flow_cnt_reg[0]  (
            .Q (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .CE (\u_touch_top/u_touch_dri/N961 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N85 ),
            .P (\u_lcd_rgb_char/u_binary2bcd_x/N0 ));
	// ../../rtl/touch/touch_dri.v:184

(* syn_encoding="onehot" *)    GTP_DFF_CE /* \u_touch_top/u_touch_dri/flow_cnt_reg[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/flow_cnt_reg[1]  (
            .Q (\u_touch_top/u_touch_dri/flow_cnt_reg [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N961 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N95 ));
	// ../../rtl/touch/touch_dri.v:184

(* syn_encoding="onehot" *)    GTP_DFF_CE /* \u_touch_top/u_touch_dri/flow_cnt_reg[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/flow_cnt_reg[2]  (
            .Q (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N961 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N102 ));
	// ../../rtl/touch/touch_dri.v:184

(* syn_encoding="onehot" *)    GTP_DFF_CE /* \u_touch_top/u_touch_dri/flow_cnt_reg[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/flow_cnt_reg[3]  (
            .Q (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N961 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N107 ));
	// ../../rtl/touch/touch_dri.v:184

(* syn_encoding="onehot" *)    GTP_DFF_CE /* \u_touch_top/u_touch_dri/flow_cnt_reg[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/flow_cnt_reg[4]  (
            .Q (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N961 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N120 ));
	// ../../rtl/touch/touch_dri.v:184

(* syn_encoding="onehot" *)    GTP_DFF_CE /* \u_touch_top/u_touch_dri/flow_cnt_reg[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/flow_cnt_reg[5]  (
            .Q (\u_touch_top/u_touch_dri/flow_cnt_reg [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N961 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N126 ));
	// ../../rtl/touch/touch_dri.v:184

(* syn_encoding="onehot" *)    GTP_DFF_CE /* \u_touch_top/u_touch_dri/flow_cnt_reg[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/flow_cnt_reg[6]  (
            .Q (\u_touch_top/u_touch_dri/flow_cnt_reg [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N961 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/_N131 ));
	// ../../rtl/touch/touch_dri.v:184

(* syn_encoding="onehot" *)    GTP_DFF_CE /* \u_touch_top/u_touch_dri/flow_cnt_reg[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/flow_cnt_reg[7]  (
            .Q (\u_touch_top/u_touch_dri/flow_cnt_reg [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N961 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N935 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/ft_flag  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/ft_flag_vname  (
            .Q (\u_touch_top/u_touch_dri/ft_flag ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (1'b1),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N11808));
    // defparam \u_touch_top/u_touch_dri/ft_flag_vname .orig_name = \u_touch_top/u_touch_dri/ft_flag ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5M /* \u_touch_top/u_touch_dri/ft_flag_ce_mux  */ #(
            .INIT(32'b00010000000000000010001000100010))
        \u_touch_top/u_touch_dri/ft_flag_ce_mux  (
            .Z (_N11808),
            .I0 (\u_touch_top/u_touch_dri/chip_version [15] ),
            .I1 (\u_touch_top/u_touch_dri/N641 ),
            .I2 (_N11956),
            .I3 (_N11960),
            .I4 (\u_touch_top/u_touch_dri/N642 ),
            .ID (\u_touch_top/u_touch_dri/ft_flag ));
	// LUT = (ID&~I1&~I4)|(~I0&~I1&I2&I3&I4) ;

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_addr[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_addr[0]  (
            .Q (\u_touch_top/i2c_addr [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1297 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1300 [0] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_addr[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_addr[1]  (
            .Q (\u_touch_top/i2c_addr [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1297 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1300 [1] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_addr[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_addr[2]  (
            .Q (\u_touch_top/i2c_addr [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1297 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1300 [2] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_addr[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_addr[3]  (
            .Q (\u_touch_top/i2c_addr [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1297 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1300 [3] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_addr[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_addr[4]  (
            .Q (\u_touch_top/i2c_addr [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1297 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1300 [4] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_addr[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_addr[5]  (
            .Q (\u_touch_top/i2c_addr [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1297 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1300 [5] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_addr[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_addr[6]  (
            .Q (\u_touch_top/i2c_addr [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1297 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1300 [6] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_addr[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_addr[7]  (
            .Q (\u_touch_top/i2c_addr [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1297 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1300 [7] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_data_w[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_data_w[1]  (
            .Q (\u_touch_top/i2c_data_w [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1216 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N933 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_data_w[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_data_w[2]  (
            .Q (\u_touch_top/i2c_data_w [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1216 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N10093));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_data_w[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_data_w[3]  (
            .Q (\u_touch_top/i2c_data_w [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1216 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N935 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT4 /* \u_touch_top/u_touch_dri/i2c_data_w[7:0]_144  */ #(
            .INIT(16'b0000000100000011))
        \u_touch_top/u_touch_dri/i2c_data_w[7:0]_144  (
            .Z (_N10093),
            .I0 (\u_touch_top/u_touch_dri/flow_cnt_reg [4] ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [2] ),
            .I2 (\u_touch_top/u_touch_dri/flow_cnt_reg [0] ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = (~I1&~I2&~I3)|(~I0&~I1&~I2) ;

    GTP_DFF_C /* \u_touch_top/u_touch_dri/i2c_exec  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_exec  (
            .Q (\u_touch_top/i2c_exec ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N394 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/i2c_rh_wl  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/i2c_rh_wl  (
            .Q (\u_touch_top/i2c_rh_wl ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1450 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1218 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/reg_num[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/reg_num[0]  (
            .Q (\u_touch_top/reg_num [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1450 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1453 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/reg_num[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/reg_num[1]  (
            .Q (\u_touch_top/reg_num [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1450 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N924 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/reg_num[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/reg_num[2]  (
            .Q (\u_touch_top/reg_num [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1450 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N945 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/slave_addr[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/slave_addr[3]  (
            .Q (\u_touch_top/slave_addr [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1074 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N9403));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/slave_addr[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/slave_addr[4]  (
            .Q (\u_touch_top/slave_addr [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1074 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (1'b1));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_C /* \u_touch_top/u_touch_dri/st_done  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/st_done_vname  (
            .Q (\u_touch_top/u_touch_dri/st_done ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N390 ));
    // defparam \u_touch_top/u_touch_dri/st_done_vname .orig_name = \u_touch_top/u_touch_dri/st_done ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/touch_int_dir  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/touch_int_dir_vname  (
            .Q (\u_touch_top/u_touch_dri/touch_int_dir ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (1'b1),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N11810));
    // defparam \u_touch_top/u_touch_dri/touch_int_dir_vname .orig_name = \u_touch_top/u_touch_dri/touch_int_dir ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT5 /* \u_touch_top/u_touch_dri/touch_int_dir_ce_mux  */ #(
            .INIT(32'b01110011011100111101000011110000))
        \u_touch_top/u_touch_dri/touch_int_dir_ce_mux  (
            .Z (_N11810),
            .I0 (\u_touch_top/u_touch_dri/N474 ),
            .I1 (\u_touch_top/u_touch_dri/st_done ),
            .I2 (\u_touch_top/u_touch_dri/touch_int_dir ),
            .I3 (\u_touch_top/u_touch_dri/cur_state_reg [1] ),
            .I4 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
	// LUT = (I1&I2&~I4)|(~I1&I4)|(~I1&I2&~I3)|(~I0&I2) ;

    GTP_LUT1 /* \u_touch_top/u_touch_dri/touch_int_dir_inv  */ #(
            .INIT(2'b01))
        \u_touch_top/u_touch_dri/touch_int_dir_inv_vname  (
            .Z (\u_touch_top/u_touch_dri/touch_int_dir_inv ),
            .I0 (\u_touch_top/u_touch_dri/touch_int_dir ));
    // defparam \u_touch_top/u_touch_dri/touch_int_dir_inv_vname .orig_name = \u_touch_top/u_touch_dri/touch_int_dir_inv ;
	// LUT = ~I0 ;

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/touch_int_out  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/touch_int_out_vname  (
            .Q (\u_touch_top/u_touch_dri/touch_int_out ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (1'b1),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N11811));
    // defparam \u_touch_top/u_touch_dri/touch_int_out_vname .orig_name = \u_touch_top/u_touch_dri/touch_int_out ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT3 /* \u_touch_top/u_touch_dri/touch_int_out_ce_mux  */ #(
            .INIT(8'b11011100))
        \u_touch_top/u_touch_dri/touch_int_out_ce_mux  (
            .Z (_N11811),
            .I0 (\u_touch_top/u_touch_dri/st_done ),
            .I1 (\u_touch_top/u_touch_dri/touch_int_out ),
            .I2 (\u_touch_top/u_touch_dri/cur_state_reg [0] ));
	// LUT = (~I0&I2)|(I1) ;

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/touch_rst_n  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/touch_rst_n  (
            .Q (nt_touch_rst_n),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N1494 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N1497 ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/touch_s_reg[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/touch_s_reg[1]  (
            .Q (\u_touch_top/u_touch_dri/touch_s_reg [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N666 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (1'b1));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/touch_valid  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/touch_valid_vname  (
            .Q (\u_touch_top/u_touch_dri/touch_valid ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (1'b1),
            .CLK (\u_touch_top/dri_clk ),
            .D (_N11809));
    // defparam \u_touch_top/u_touch_dri/touch_valid_vname .orig_name = \u_touch_top/u_touch_dri/touch_valid ;
	// ../../rtl/touch/touch_dri.v:184

    GTP_LUT4 /* \u_touch_top/u_touch_dri/touch_valid_ce_mux  */ #(
            .INIT(16'b1011100011110000))
        \u_touch_top/u_touch_dri/touch_valid_ce_mux  (
            .Z (_N11809),
            .I0 (\u_touch_top/u_touch_dri/N296 ),
            .I1 (\u_touch_top/u_touch_dri/flow_cnt_reg [3] ),
            .I2 (\u_touch_top/u_touch_dri/touch_valid ),
            .I3 (\u_touch_top/u_touch_dri/next_state [4] ));
	// LUT = (I2&~I3)|(I0&I1&I3)|(~I1&I2) ;

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[0]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [0] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[1]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [1] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[2]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [2] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[3]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [3] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[4]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [4] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[5]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [5] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[6]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [6] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[7]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [7] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[8]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [8] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[9]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [9] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[10]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [10] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[11]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [11] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[12]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [12] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [12] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[13]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [13] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [13] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[14]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [14] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [14] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord[15]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord [15] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N376 [15] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[0]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N716 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [0] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[1]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N716 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [1] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[2]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N716 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [2] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[3]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N716 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [3] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[4]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N716 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [4] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[5]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N716 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [5] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[6]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N716 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [6] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[7]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N716 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [7] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[8]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N739 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [0] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[9]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N739 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [1] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[10]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N739 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [2] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[11]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N739 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [3] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[12]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [12] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N739 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [4] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[13]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [13] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N739 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [5] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[14]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [14] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N739 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [6] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_x_coord_t[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_x_coord_t[15]  (
            .Q (\u_touch_top/u_touch_dri/tp_x_coord_t [15] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N739 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [7] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[0]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [0] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[1]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [1] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[2]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [2] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[3]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [3] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[4]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [4] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[5]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [5] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[6]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [6] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[7]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [7] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[8]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [8] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[9]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [9] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[10]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [10] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[11]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [11] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[12]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [12] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [12] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[13]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [13] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [13] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[14]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [14] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [14] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord[15]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord [15] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/next_state [6] ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/u_touch_dri/N377 [15] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[0]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[0]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [0] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N948 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [0] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[1]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[1]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [1] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N948 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [1] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[2]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[2]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [2] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N948 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [2] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[3]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[3]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [3] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N948 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [3] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[4]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[4]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [4] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N948 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [4] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[5]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[5]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [5] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N948 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [5] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[6]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[6]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [6] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N948 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [6] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[7]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[7]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [7] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N948 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [7] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[8]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[8]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [8] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N614 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [0] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[9]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[9]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [9] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N614 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [1] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[10]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[10]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [10] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N614 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [2] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[11]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[11]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [11] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N614 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [3] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[12]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[12]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [12] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N614 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [4] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[13]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[13]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [13] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N614 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [5] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[14]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[14]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [14] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N614 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [6] ));
	// ../../rtl/touch/touch_dri.v:184

    GTP_DFF_CE /* \u_touch_top/u_touch_dri/tp_y_coord_t[15]  */ #(
            .GRS_EN("TRUE"), 
            .INIT(1'b0))
        \u_touch_top/u_touch_dri/tp_y_coord_t[15]  (
            .Q (\u_touch_top/u_touch_dri/tp_y_coord_t [15] ),
            .C (\u_lcd_rgb_char/u_binary2bcd_x/N0 ),
            .CE (\u_touch_top/u_touch_dri/N614 ),
            .CLK (\u_touch_top/dri_clk ),
            .D (\u_touch_top/i2c_data_r [7] ));
	// ../../rtl/touch/touch_dri.v:184


endmodule

