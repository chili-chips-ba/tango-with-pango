//****************************************Copyright (c)***********************************//
//ԭ�Ӹ����߽�ѧƽ̨��www.yuanzige.com
//����֧�֣�http://www.openedv.com/forum.php
//�Ա����̣�https://zhengdianyuanzi.tmall.com
//��ע΢�Ź���ƽ̨΢�źţ�"����ԭ��"����ѻ�ȡZYNQ & FPGA & STM32 & LINUX���ϡ�
//��Ȩ���У�����ؾ���
//Copyright(C) ����ԭ�� 2023-2033
//All rights reserved                                  
//----------------------------------------------------------------------------------------
// File name:           tb_led
// Created by:          ����ԭ��
// Created date:        2023��3��30��11:12:36
// Version:             V1.0
// Descriptions:        ����LEDʵ�鼤���ļ�
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

`timescale 1ns / 1ns        //���浥λ/���澫��

module tb_led();

//reg define
reg           key;
//wire define
wire          led;

//�źų�ʼ��
initial begin
    key <= 1'b1;   //�����ϵ�Ĭ�ϸߵ�ƽ

//key�źű仯
    #200           //�ӳ�200ns
    key <= 1'b1;   //����û�б�����
    #1000  
    key <= 1'b0;   //����������
    #600  
    key <= 1'b1;
    #1000  
    key <= 1'b0;
end

//����ledģ��
led  u_led(
    .key          (key),
    .led          (led)
    );

endmodule

