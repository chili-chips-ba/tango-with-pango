//****************************************Copyright (c)***********************************//
//ԭ�Ӹ����߽�ѧƽ̨��www.yuanzige.com
//����֧�֣�http://www.openedv.com/forum.php
//�Ա����̣�https://zhengdianyuanzi.tmall.com
//��ע΢�Ź���ƽ̨΢�źţ�"����ԭ��"����ѻ�ȡZYNQ & FPGA & STM32 & LINUX���ϡ�
//��Ȩ���У�����ؾ���
//Copyright(C) ����ԭ�� 2023-2033
//All rights reserved                                  
//----------------------------------------------------------------------------------------
// File name:           led
// Created by:          ����ԭ��
// Created date:        2023��3��30��09:40:02
// Version:             V1.0
// Descriptions:        ����LED��ʵ��
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module led(                     
    input     key , //���밴��
    
    output    led   //���led��
);

//*****************************************************
//**                  main code
//*****************************************************

//�ϵ簴��Ĭ�ϸߵ�ƽ��led�Ʊ��ֳ���
//���������£�����ֵΪ�͵�ƽ��led�Ʊ�����
assign led = ~key;    //��������ֵȡ����ֵ��led��

endmodule